// Fix_Add.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module Fix_Add (
		input  wire        clk,    //    clk.clk
		input  wire        rst,    //    rst.reset
		input  wire [0:0]  en,     //     en.en
		input  wire [31:0] a0,     //     a0.a0
		input  wire [31:0] a1,     //     a1.a1
		output wire [32:0] result  // result.result
	);

	Fix_Add_altera_fxp_functions_191_i22v3ci fxp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.rst    (rst),    //   input,   width = 1,    rst.reset
		.en     (en),     //   input,   width = 1,     en.en
		.a0     (a0),     //   input,  width = 32,     a0.a0
		.a1     (a1),     //   input,  width = 32,     a1.a1
		.result (result)  //  output,  width = 33, result.result
	);

endmodule
