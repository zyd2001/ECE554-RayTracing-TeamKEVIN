// Fix_Mul.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module Fix_Mul (
		input  wire        clk,    //    clk.clk
		input  wire        rst,    //    rst.reset
		input  wire [0:0]  en,     //     en.en
		input  wire [31:0] a,      //      a.a
		input  wire [31:0] b,      //      b.b
		output wire [63:0] result  // result.result
	);

	Fix_Mul_altera_fxp_functions_191_vsvne7a fxp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.rst    (rst),    //   input,   width = 1,    rst.reset
		.en     (en),     //   input,   width = 1,     en.en
		.a      (a),      //   input,  width = 32,      a.a
		.b      (b),      //   input,  width = 32,      b.b
		.result (result)  //  output,  width = 64, result.result
	);

endmodule
