module Fix_Add (
		input  wire        clk,    //    clk.clk
		input  wire        rst,    //    rst.reset
		input  wire [0:0]  en,     //     en.en
		input  wire [31:0] a0,     //     a0.a0
		input  wire [31:0] a1,     //     a1.a1
		output wire [32:0] result  // result.result
	);
endmodule

