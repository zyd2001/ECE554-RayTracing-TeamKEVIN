module Fix_Sqrt (
		input  wire        clk,     //     clk.clk
		input  wire        rst,     //     rst.reset
		input  wire [0:0]  en,      //      en.en
		input  wire [31:0] radical, // radical.radical
		output wire [31:0] result   //  result.result
	);
endmodule

