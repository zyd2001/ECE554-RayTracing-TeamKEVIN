// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/20/2021 23:05:55"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Float_Sqrt (
	q,
	clk,
	areset,
	en,
	a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	clk;
input 	areset;
input 	[0:0] en;
input 	[31:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a8_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a9_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a10_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a11_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a12_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a13_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a14_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a15_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a16_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a17_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a18_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a19_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a20_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a21_a_aq;
wire fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a22_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aadd_7_a1_sumout;
wire fp_functions_0_aadd_7_a2;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a1_a_aq;
wire fp_functions_0_aadd_7_a6_sumout;
wire fp_functions_0_aadd_7_a7;
wire fp_functions_0_aadd_7_a11_sumout;
wire fp_functions_0_aadd_7_a12;
wire fp_functions_0_aadd_7_a16_sumout;
wire fp_functions_0_aadd_7_a17;
wire fp_functions_0_aadd_7_a21_sumout;
wire fp_functions_0_aadd_7_a22;
wire fp_functions_0_aadd_7_a26_sumout;
wire fp_functions_0_aadd_7_a27;
wire fp_functions_0_aadd_7_a31_sumout;
wire fp_functions_0_aadd_7_a32;
wire fp_functions_0_aadd_7_a36_sumout;
wire fp_functions_0_aadd_7_a37;
wire fp_functions_0_aadd_7_a41_sumout;
wire fp_functions_0_aadd_7_a42;
wire fp_functions_0_aadd_7_a46_sumout;
wire fp_functions_0_aadd_7_a47;
wire fp_functions_0_aadd_7_a51_sumout;
wire fp_functions_0_aadd_7_a52;
wire fp_functions_0_aadd_7_a56_sumout;
wire fp_functions_0_aadd_7_a57;
wire fp_functions_0_aadd_7_a61_sumout;
wire fp_functions_0_aadd_7_a62;
wire fp_functions_0_aadd_7_a66_sumout;
wire fp_functions_0_aadd_7_a67;
wire fp_functions_0_aadd_7_a71_sumout;
wire fp_functions_0_aadd_7_a72;
wire fp_functions_0_aadd_7_a76_sumout;
wire fp_functions_0_aadd_7_a77;
wire fp_functions_0_aadd_7_a81_sumout;
wire fp_functions_0_aadd_7_a82;
wire fp_functions_0_aadd_7_a86_sumout;
wire fp_functions_0_aadd_7_a87;
wire fp_functions_0_aadd_7_a91_sumout;
wire fp_functions_0_aadd_7_a92;
wire fp_functions_0_aadd_7_a96_sumout;
wire fp_functions_0_aadd_7_a97;
wire fp_functions_0_aadd_7_a101_sumout;
wire fp_functions_0_aadd_7_a102;
wire fp_functions_0_aadd_7_a106_sumout;
wire fp_functions_0_aadd_7_a107;
wire fp_functions_0_aadd_7_a111_sumout;
wire fp_functions_0_aadd_7_a112;
wire fp_functions_0_aadd_12_a1_sumout;
wire fp_functions_0_aadd_12_a2;
wire fp_functions_0_aadd_12_a6_sumout;
wire fp_functions_0_aadd_12_a7;
wire fp_functions_0_aadd_12_a11_sumout;
wire fp_functions_0_aadd_12_a12;
wire fp_functions_0_aadd_12_a16_sumout;
wire fp_functions_0_aadd_12_a17;
wire fp_functions_0_aadd_12_a21_sumout;
wire fp_functions_0_aadd_12_a22;
wire fp_functions_0_aadd_12_a26_sumout;
wire fp_functions_0_aadd_12_a27;
wire fp_functions_0_aadd_12_a31_sumout;
wire fp_functions_0_aadd_12_a32;
wire fp_functions_0_aadd_12_a36_sumout;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_aadd_7_a117_cout;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a1_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a;
wire fp_functions_0_aadd_7_a121_sumout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a24_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a25_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a26_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a27_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a28_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a29_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a30_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a31_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a32_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a33_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a34_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a35_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a36_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a37_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a38_a;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_aadd_7_a127_cout;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a1_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a;
wire fp_functions_0_aadd_7_a132_cout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_aadd_7_a137_cout;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a1_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist1_lowRangeB_uid76_invPolyEval_b_1_q_a0_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a0_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a1_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a2_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a3_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a4_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a5_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a6_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a7_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a8_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a9_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a10_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a11_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a12_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a13_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a14_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a15_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a16_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a17_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a18_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a19_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a20_a_aq;
wire fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a21_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a8_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a9_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a10_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a11_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a12_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a13_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a14_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a15_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_aadd_7_a142_cout;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a0_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a1_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a2_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a3_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a4_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a5_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a6_a_aq;
wire fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a7_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aadd_2_a1_sumout;
wire fp_functions_0_aadd_2_a2;
wire fp_functions_0_aadd_2_a6_sumout;
wire fp_functions_0_aadd_2_a7;
wire fp_functions_0_aadd_2_a11_sumout;
wire fp_functions_0_aadd_2_a12;
wire fp_functions_0_aadd_2_a16_sumout;
wire fp_functions_0_aadd_2_a17;
wire fp_functions_0_aadd_2_a21_sumout;
wire fp_functions_0_aadd_2_a22;
wire fp_functions_0_aadd_2_a26_sumout;
wire fp_functions_0_aadd_2_a27;
wire fp_functions_0_aadd_2_a31_sumout;
wire fp_functions_0_aadd_2_a32;
wire fp_functions_0_aadd_2_a36_sumout;
wire fp_functions_0_aadd_2_a37;
wire fp_functions_0_aadd_2_a41_sumout;
wire fp_functions_0_aadd_2_a42;
wire fp_functions_0_aadd_2_a46_sumout;
wire fp_functions_0_aadd_2_a47;
wire fp_functions_0_aadd_2_a51_sumout;
wire fp_functions_0_aadd_2_a52;
wire fp_functions_0_aadd_2_a56_sumout;
wire fp_functions_0_aadd_2_a57;
wire fp_functions_0_aadd_2_a61_sumout;
wire fp_functions_0_aadd_2_a62;
wire fp_functions_0_aadd_2_a66_sumout;
wire fp_functions_0_aadd_2_a67;
wire fp_functions_0_aadd_2_a71_sumout;
wire fp_functions_0_aadd_2_a72;
wire fp_functions_0_aadd_2_a76_sumout;
wire fp_functions_0_aadd_2_a77;
wire fp_functions_0_aadd_2_a81_sumout;
wire fp_functions_0_aadd_2_a82;
wire fp_functions_0_aadd_2_a86_sumout;
wire fp_functions_0_aadd_2_a87;
wire fp_functions_0_aadd_2_a91_sumout;
wire fp_functions_0_aadd_2_a92;
wire fp_functions_0_aadd_2_a96_sumout;
wire fp_functions_0_aadd_2_a97;
wire fp_functions_0_aadd_2_a101_sumout;
wire fp_functions_0_aadd_2_a102;
wire fp_functions_0_aadd_2_a106_sumout;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_cmpReg_q_a0_a_aq;
wire fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq_aq;
wire fp_functions_0_aadd_10_a1_sumout;
wire fp_functions_0_aadd_10_a2;
wire fp_functions_0_aadd_10_a6_sumout;
wire fp_functions_0_aadd_10_a7;
wire fp_functions_0_aadd_10_a11_sumout;
wire fp_functions_0_aadd_10_a12;
wire fp_functions_0_aadd_10_a16_sumout;
wire fp_functions_0_aadd_10_a17;
wire fp_functions_0_aadd_10_a21_sumout;
wire fp_functions_0_aadd_10_a22;
wire fp_functions_0_aadd_10_a26_sumout;
wire fp_functions_0_aadd_10_a27;
wire fp_functions_0_aadd_10_a31_sumout;
wire fp_functions_0_aadd_10_a32;
wire fp_functions_0_aadd_10_a36_sumout;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA24;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA25;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA26;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA27;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA28;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA29;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA30;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA31;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA32;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA33;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA34;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA35;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA36;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a1_a_aq;
wire fp_functions_0_aadd_10_a42_cout;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a0_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a1_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a2_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a3_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a4_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a5_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a6_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a7_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a8_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a9_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a10_a_aq;
wire fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a11_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a0_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a1_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a2_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a3_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a4_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a5_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a6_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a7_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a8_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a9_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a10_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a11_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a12_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a13_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a14_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a15_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a0_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a1_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a2_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a3_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a4_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a5_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a6_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a7_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a8_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a9_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a10_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a11_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a12_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a13_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a14_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a15_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a0_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a1_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a2_a_aq;
wire fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a3_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a1_a_aq;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_afracSel_uid48_fpSqrtTest_q_a1_a_aq;
wire fp_functions_0_anegZero_uid59_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_afracXIsZero_uid15_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a_aq;
wire fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aMux_32_a2_combout;
wire fp_functions_0_aMux_31_a0_combout;
wire fp_functions_0_aMux_30_a0_combout;
wire fp_functions_0_aMux_29_a0_combout;
wire fp_functions_0_aMux_28_a0_combout;
wire fp_functions_0_aMux_27_a0_combout;
wire fp_functions_0_aMux_26_a0_combout;
wire fp_functions_0_aMux_25_a0_combout;
wire fp_functions_0_aMux_24_a0_combout;
wire fp_functions_0_aMux_23_a0_combout;
wire fp_functions_0_aMux_22_a0_combout;
wire fp_functions_0_aMux_21_a0_combout;
wire fp_functions_0_aMux_20_a0_combout;
wire fp_functions_0_aMux_19_a0_combout;
wire fp_functions_0_aMux_18_a0_combout;
wire fp_functions_0_aMux_17_a0_combout;
wire fp_functions_0_aMux_16_a0_combout;
wire fp_functions_0_aMux_15_a0_combout;
wire fp_functions_0_aMux_14_a0_combout;
wire fp_functions_0_aMux_13_a0_combout;
wire fp_functions_0_aMux_12_a0_combout;
wire fp_functions_0_aMux_11_a0_combout;
wire fp_functions_0_aMux_10_a0_combout;
wire fp_functions_0_aMux_9_a2_combout;
wire fp_functions_0_aMux_9_a3_combout;
wire fp_functions_0_aMux_9_a4_combout;
wire fp_functions_0_aMux_9_a5_combout;
wire fp_functions_0_aMux_9_a6_combout;
wire fp_functions_0_aMux_9_a7_combout;
wire fp_functions_0_aMux_9_a8_combout;
wire fp_functions_0_aMux_9_a9_combout;
wire fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq;
wire fp_functions_0_ai1410_a0_combout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fp_functions_0_ai1568_a0_combout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0_combout;
wire fp_functions_0_ai1568_a1_combout;
wire fp_functions_0_ai1568_a2_combout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1_combout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2_combout;
wire fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3_combout;
wire fp_functions_0_areduce_nor_11_acombout;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai1109_a0_combout;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fp_functions_0_ai1424_a0_combout;
wire fp_functions_0_aadd_8_a0_combout;
wire fp_functions_0_aadd_8_a1_combout;
wire fp_functions_0_aadd_8_a2_combout;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai1140_a0_combout;
wire fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_5_acombout;
wire fp_functions_0_areduce_nor_8_acombout;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai768_a0_combout;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq;
wire fp_functions_0_ai1121_a0_combout;
wire fp_functions_0_ai1121_a1_combout;
wire fp_functions_0_ai1121_a2_combout;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai799_a0_combout;
wire fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_3_acombout;
wire fp_functions_0_areduce_nor_6_acombout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout;
wire fp_functions_0_ai780_a0_combout;
wire fp_functions_0_ai780_a1_combout;
wire fp_functions_0_ai780_a2_combout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai481_a0_combout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_areduce_nor_4_acombout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai513_a0_combout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_1_acombout;
wire fp_functions_0_ai493_a0_combout;
wire fp_functions_0_ai493_a1_combout;
wire fp_functions_0_ai493_a2_combout;
wire fp_functions_0_areduce_nor_2_acombout;
wire fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a_aq;
wire fp_functions_0_aMux_1_a0_combout;
wire fp_functions_0_ai1741_a0_combout;
wire fp_functions_0_aMux_1_a1_combout;
wire fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a_acombout;
wire fp_functions_0_areduce_nor_9_a0_combout;
wire fp_functions_0_areduce_nor_9_acombout;
wire fp_functions_0_areduce_nor_10_a0_combout;
wire fp_functions_0_areduce_nor_10_a1_combout;
wire fp_functions_0_areduce_nor_10_a2_combout;
wire fp_functions_0_areduce_nor_10_a3_combout;
wire fp_functions_0_areduce_nor_10_acombout;
wire fp_functions_0_areduce_nor_0_a0_combout;
wire fp_functions_0_areduce_nor_0_acombout;
wire fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0_combout;
wire a_a23_a_a_wirecell_combout;

wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus;
wire [63:0] fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [63:0] fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus[0];

assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a0_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a1_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a2_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a3_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a4_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a5_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a6_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a7_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a8_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a9_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a10_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a11_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a12_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a13_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a14_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a15_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a16_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a17_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a18_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a19_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a20_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a21_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a22_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a23_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a24_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a25_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a26_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a27_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a28_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a29_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a30_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a31_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a32_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a33_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a34_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a35_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a36_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a37_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a38_a = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA39 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA40 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA41 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA42 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA43 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA44 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA45 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA46 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA47 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA48 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA49 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a0_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a1_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a2_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a3_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a4_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a5_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a6_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a7_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a8_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a9_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a10_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a11_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a12_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a13_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a14_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a15_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a16_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a17_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a18_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a19_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a20_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a21_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a22_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a23_a = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA24 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA25 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA26 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA27 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA28 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA29 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA30 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA31 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA32 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA33 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA34 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA35 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA36 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA37 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA38 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA39 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA40 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA41 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA42 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA43 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA44 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA45 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA46 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA47 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA48 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA49 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19 = fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_7_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_12_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_7_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a117_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a1_sumout),
	.cout(fp_functions_0_aadd_7_a2),
	.shareout());
defparam fp_functions_0_aadd_7_a1.extended_lut = "off";
defparam fp_functions_0_aadd_7_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a1.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a1_a_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_7_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a6_sumout),
	.cout(fp_functions_0_aadd_7_a7),
	.shareout());
defparam fp_functions_0_aadd_7_a6.extended_lut = "off";
defparam fp_functions_0_aadd_7_a6.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a11_sumout),
	.cout(fp_functions_0_aadd_7_a12),
	.shareout());
defparam fp_functions_0_aadd_7_a11.extended_lut = "off";
defparam fp_functions_0_aadd_7_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a16_sumout),
	.cout(fp_functions_0_aadd_7_a17),
	.shareout());
defparam fp_functions_0_aadd_7_a16.extended_lut = "off";
defparam fp_functions_0_aadd_7_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a21_sumout),
	.cout(fp_functions_0_aadd_7_a22),
	.shareout());
defparam fp_functions_0_aadd_7_a21.extended_lut = "off";
defparam fp_functions_0_aadd_7_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a26_sumout),
	.cout(fp_functions_0_aadd_7_a27),
	.shareout());
defparam fp_functions_0_aadd_7_a26.extended_lut = "off";
defparam fp_functions_0_aadd_7_a26.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a31_sumout),
	.cout(fp_functions_0_aadd_7_a32),
	.shareout());
defparam fp_functions_0_aadd_7_a31.extended_lut = "off";
defparam fp_functions_0_aadd_7_a31.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a36_sumout),
	.cout(fp_functions_0_aadd_7_a37),
	.shareout());
defparam fp_functions_0_aadd_7_a36.extended_lut = "off";
defparam fp_functions_0_aadd_7_a36.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a41_sumout),
	.cout(fp_functions_0_aadd_7_a42),
	.shareout());
defparam fp_functions_0_aadd_7_a41.extended_lut = "off";
defparam fp_functions_0_aadd_7_a41.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a46_sumout),
	.cout(fp_functions_0_aadd_7_a47),
	.shareout());
defparam fp_functions_0_aadd_7_a46.extended_lut = "off";
defparam fp_functions_0_aadd_7_a46.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a51_sumout),
	.cout(fp_functions_0_aadd_7_a52),
	.shareout());
defparam fp_functions_0_aadd_7_a51.extended_lut = "off";
defparam fp_functions_0_aadd_7_a51.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a56_sumout),
	.cout(fp_functions_0_aadd_7_a57),
	.shareout());
defparam fp_functions_0_aadd_7_a56.extended_lut = "off";
defparam fp_functions_0_aadd_7_a56.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a61_sumout),
	.cout(fp_functions_0_aadd_7_a62),
	.shareout());
defparam fp_functions_0_aadd_7_a61.extended_lut = "off";
defparam fp_functions_0_aadd_7_a61.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a66_sumout),
	.cout(fp_functions_0_aadd_7_a67),
	.shareout());
defparam fp_functions_0_aadd_7_a66.extended_lut = "off";
defparam fp_functions_0_aadd_7_a66.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a71_sumout),
	.cout(fp_functions_0_aadd_7_a72),
	.shareout());
defparam fp_functions_0_aadd_7_a71.extended_lut = "off";
defparam fp_functions_0_aadd_7_a71.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a76_sumout),
	.cout(fp_functions_0_aadd_7_a77),
	.shareout());
defparam fp_functions_0_aadd_7_a76.extended_lut = "off";
defparam fp_functions_0_aadd_7_a76.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a81_sumout),
	.cout(fp_functions_0_aadd_7_a82),
	.shareout());
defparam fp_functions_0_aadd_7_a81.extended_lut = "off";
defparam fp_functions_0_aadd_7_a81.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a86_sumout),
	.cout(fp_functions_0_aadd_7_a87),
	.shareout());
defparam fp_functions_0_aadd_7_a86.extended_lut = "off";
defparam fp_functions_0_aadd_7_a86.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a91(
	.dataa(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a91_sumout),
	.cout(fp_functions_0_aadd_7_a92),
	.shareout());
defparam fp_functions_0_aadd_7_a91.extended_lut = "off";
defparam fp_functions_0_aadd_7_a91.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_7_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a96(
	.dataa(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a96_sumout),
	.cout(fp_functions_0_aadd_7_a97),
	.shareout());
defparam fp_functions_0_aadd_7_a96.extended_lut = "off";
defparam fp_functions_0_aadd_7_a96.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_7_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a101(
	.dataa(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a101_sumout),
	.cout(fp_functions_0_aadd_7_a102),
	.shareout());
defparam fp_functions_0_aadd_7_a101.extended_lut = "off";
defparam fp_functions_0_aadd_7_a101.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_7_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a106(
	.dataa(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a106_sumout),
	.cout(fp_functions_0_aadd_7_a107),
	.shareout());
defparam fp_functions_0_aadd_7_a106.extended_lut = "off";
defparam fp_functions_0_aadd_7_a106.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_7_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a111(
	.dataa(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a111_sumout),
	.cout(fp_functions_0_aadd_7_a112),
	.shareout());
defparam fp_functions_0_aadd_7_a111.extended_lut = "off";
defparam fp_functions_0_aadd_7_a111.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_7_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_7_a121_sumout),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a1_sumout),
	.cout(fp_functions_0_aadd_12_a2),
	.shareout());
defparam fp_functions_0_aadd_12_a1.extended_lut = "off";
defparam fp_functions_0_aadd_12_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_12_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a6_sumout),
	.cout(fp_functions_0_aadd_12_a7),
	.shareout());
defparam fp_functions_0_aadd_12_a6.extended_lut = "off";
defparam fp_functions_0_aadd_12_a6.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a11_sumout),
	.cout(fp_functions_0_aadd_12_a12),
	.shareout());
defparam fp_functions_0_aadd_12_a11.extended_lut = "off";
defparam fp_functions_0_aadd_12_a11.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a16_sumout),
	.cout(fp_functions_0_aadd_12_a17),
	.shareout());
defparam fp_functions_0_aadd_12_a16.extended_lut = "off";
defparam fp_functions_0_aadd_12_a16.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a21_sumout),
	.cout(fp_functions_0_aadd_12_a22),
	.shareout());
defparam fp_functions_0_aadd_12_a21.extended_lut = "off";
defparam fp_functions_0_aadd_12_a21.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a26_sumout),
	.cout(fp_functions_0_aadd_12_a27),
	.shareout());
defparam fp_functions_0_aadd_12_a26.extended_lut = "off";
defparam fp_functions_0_aadd_12_a26.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a31_sumout),
	.cout(fp_functions_0_aadd_12_a32),
	.shareout());
defparam fp_functions_0_aadd_12_a31.extended_lut = "off";
defparam fp_functions_0_aadd_12_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_12_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_12_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_12_a36_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_12_a36.extended_lut = "off";
defparam fp_functions_0_aadd_12_a36.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_12_a36.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "01B24401E772568BE9BDD8700362DF596AA0DDE9CF8B22F29F710E916D060190";

fourteennm_lcell_comb fp_functions_0_aadd_7_a117(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a127_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_7_a117_cout),
	.shareout());
defparam fp_functions_0_aadd_7_a117.extended_lut = "off";
defparam fp_functions_0_aadd_7_a117.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a117.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a2_a_a1_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "272D7B7CE4AF822F54384D2F1C923607E8C9B6809CFDBC68C92DD158EAEBC7BC";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "310728184CAEB84D5C0F8CD074FA301E36596BEFBE326A546C86136332672E78";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "3B242B702317E42485BAB58AEAFEE58ABE39A229E6E14CC4E8E8181B43061F30";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "3D993AB9864917E3ED5FE1ACA29A469FF2CAFAF5BCEA7093537CD1D983A599E0";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "94819B7C25B6C1866E8EE99A63944BF11F2912433DB380E53D0B590130FF0F40";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "BF4D1DCDAA492243CD04E4D3499A6239927B91190F5A669FCD6B45701EE8AF2A";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "FBB596E0171C724DBF9BD085EB50104F665A98432114F06EE0AFD0B93829FC2A";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "D7D230A17AEBACCBDE9744C45058EDB651919D3D9E4F50A0A16D24298239746E";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "E54FDA61A9F29F67EA6539B93D220BD0CFE2CB01D53F9A60CB11AC337C99AC46";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "F99549E1CD567F8AA606547E54FCA7E56AA9B8FE19AAB61F0DAB63C2558636DE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "FE1992B4A4CE000CCB52CC0066AA6006D99878001E3324AAA498E003992A923E";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "FFE1E3393694AAA5A6CE3C0078CCB552387807FFE03C38CCC92D4AA94B6671FE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "FFFE03C1C718CCC93494A9552A5A6CCEAD52AAAAAA956A5A5B64D998C71E0FFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "FFFFFC01F81F0F0E38E73199B36CB69464C99999998CE639C71C38783F01FFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "55555554AAB55AA56A5294B496DA6DB2B692D2D2D2D6B4AD6A56AD52AA555554";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "9999999933266CC9B364D926DB6CB6DB38E31CE31CE738CE7398CE6333999998";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_bit_number = 21;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_bit_number = 21;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mem_init0 = "E1E1E1E1C3C78F0E3C78E1C71C70C71C3F03E0FC1F07C0F07C1F0F83C3E1E1E0";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_bit_number = 22;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_bit_number = 22;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mem_init0 = "FE01FE01FC07F00FC07F01F81F80F81FC003FF001FF800FF801FF003FC01FE00";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_bit_number = 23;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_bit_number = 23;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mem_init0 = "FFFE0001FFF8000FFF8001FFE000FFE00003FFFFE00000FFFFE00003FFFE0000";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_bit_number = 24;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_bit_number = 24;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mem_init0 = "FFFFFFFE0000000FFFFFFE000000FFFFFFFC0000000000FFFFFFFFFC00000000";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_bit_number = 25;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_bit_number = 25;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mem_init0 = "FFFFFFFFFFFFFFF0000000000000FFFFFFFFFFFFFFFFFF000000000000000000";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_bit_number = 26;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_bit_number = 26;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000";

fourteennm_lcell_comb fp_functions_0_aadd_7_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a132_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a121_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_7_a121.extended_lut = "off";
defparam fp_functions_0_aadd_7_a121.lut_mask = 64'h0000000000000FF0;
defparam fp_functions_0_aadd_7_a121.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a22_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a21_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a20_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a19_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a18_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a17_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a16_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a15_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a14_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a13_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a12_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a11_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a10_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a8_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a7_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a5_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a4_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a2_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a1_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a15_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a14_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a13_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a12_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout,fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout,
fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.ax_width = 23;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.ay_scan_in_width = 16;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.operation_mode = "m27x27";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.result_a_width = 39;
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.signed_max = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "BF8E327A079B0D5B0CB27788D52FE2B35A79C681C1F69E695978A238D34DF67A";

fourteennm_lcell_comb fp_functions_0_aadd_7_a127(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a137_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_7_a127_cout),
	.shareout());
defparam fp_functions_0_aadd_7_a127.extended_lut = "off";
defparam fp_functions_0_aadd_7_a127.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a127.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a3_a_a1_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_bit_number = 28;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_bit_number = 28;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

fourteennm_lcell_comb fp_functions_0_aadd_7_a132(
	.dataa(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a112),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_7_a132_cout),
	.shareout());
defparam fp_functions_0_aadd_7_a132.extended_lut = "off";
defparam fp_functions_0_aadd_7_a132.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_7_a132.shared_arith = "off";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1410_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 4;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 13;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 14;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist10_exprmux_uid31_fpsqrttest_q_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "27D4297CA8AE58C351BE55DB8A688E6D8FBF4D3A6257DB6153EC267435E8A37D";

fourteennm_lcell_comb fp_functions_0_aadd_7_a137(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a142_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_7_a137_cout),
	.shareout());
defparam fp_functions_0_aadd_7_a137.extended_lut = "off";
defparam fp_functions_0_aadd_7_a137.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a137.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a4_a_a1_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_bit_number = 27;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_bit_number = 27;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_11_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_lowRangeB_uid76_invPolyEval_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_lowRangeB_uid76_invPolyEval_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist1_lowRangeB_uid76_invPolyEval_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_lowRangeB_uid76_invPolyEval_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a0_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a1_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a2_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a3_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a4_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a5_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a6_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a7_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a8_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a9_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a10_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a11_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a12_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a13_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a14_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a15_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a16_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a17_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a18_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a19_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a20_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a21_a_aq));
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a8_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a9_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a10_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a11_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a12_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a13_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a14_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a15_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a15_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1109_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist9_yaddr_uid35_fpsqrttest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "09CCF058A4275C06A943D5272B9A66AC73E857E05BBCE62D49160A014123EF98";

fourteennm_lcell_comb fp_functions_0_aadd_7_a142(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_7_a142_cout),
	.shareout());
defparam fp_functions_0_aadd_7_a142.extended_lut = "off";
defparam fp_functions_0_aadd_7_a142.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a142.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a5_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1424_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_8_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_8_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_8_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a0_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a1_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a2_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a3_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a4_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a5_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a6_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_10_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a7_a_aq));
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a1_sumout),
	.cout(fp_functions_0_aadd_2_a2),
	.shareout());
defparam fp_functions_0_aadd_2_a1.extended_lut = "off";
defparam fp_functions_0_aadd_2_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a6_sumout),
	.cout(fp_functions_0_aadd_2_a7),
	.shareout());
defparam fp_functions_0_aadd_2_a6.extended_lut = "off";
defparam fp_functions_0_aadd_2_a6.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a11_sumout),
	.cout(fp_functions_0_aadd_2_a12),
	.shareout());
defparam fp_functions_0_aadd_2_a11.extended_lut = "off";
defparam fp_functions_0_aadd_2_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a16_sumout),
	.cout(fp_functions_0_aadd_2_a17),
	.shareout());
defparam fp_functions_0_aadd_2_a16.extended_lut = "off";
defparam fp_functions_0_aadd_2_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a21_sumout),
	.cout(fp_functions_0_aadd_2_a22),
	.shareout());
defparam fp_functions_0_aadd_2_a21.extended_lut = "off";
defparam fp_functions_0_aadd_2_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a26_sumout),
	.cout(fp_functions_0_aadd_2_a27),
	.shareout());
defparam fp_functions_0_aadd_2_a26.extended_lut = "off";
defparam fp_functions_0_aadd_2_a26.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a31_sumout),
	.cout(fp_functions_0_aadd_2_a32),
	.shareout());
defparam fp_functions_0_aadd_2_a31.extended_lut = "off";
defparam fp_functions_0_aadd_2_a31.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a36_sumout),
	.cout(fp_functions_0_aadd_2_a37),
	.shareout());
defparam fp_functions_0_aadd_2_a36.extended_lut = "off";
defparam fp_functions_0_aadd_2_a36.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a41_sumout),
	.cout(fp_functions_0_aadd_2_a42),
	.shareout());
defparam fp_functions_0_aadd_2_a41.extended_lut = "off";
defparam fp_functions_0_aadd_2_a41.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a46_sumout),
	.cout(fp_functions_0_aadd_2_a47),
	.shareout());
defparam fp_functions_0_aadd_2_a46.extended_lut = "off";
defparam fp_functions_0_aadd_2_a46.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a51_sumout),
	.cout(fp_functions_0_aadd_2_a52),
	.shareout());
defparam fp_functions_0_aadd_2_a51.extended_lut = "off";
defparam fp_functions_0_aadd_2_a51.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a56_sumout),
	.cout(fp_functions_0_aadd_2_a57),
	.shareout());
defparam fp_functions_0_aadd_2_a56.extended_lut = "off";
defparam fp_functions_0_aadd_2_a56.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_2_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a61(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a61_sumout),
	.cout(fp_functions_0_aadd_2_a62),
	.shareout());
defparam fp_functions_0_aadd_2_a61.extended_lut = "off";
defparam fp_functions_0_aadd_2_a61.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a66(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a66_sumout),
	.cout(fp_functions_0_aadd_2_a67),
	.shareout());
defparam fp_functions_0_aadd_2_a66.extended_lut = "off";
defparam fp_functions_0_aadd_2_a66.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a71(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a71_sumout),
	.cout(fp_functions_0_aadd_2_a72),
	.shareout());
defparam fp_functions_0_aadd_2_a71.extended_lut = "off";
defparam fp_functions_0_aadd_2_a71.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a76(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a76_sumout),
	.cout(fp_functions_0_aadd_2_a77),
	.shareout());
defparam fp_functions_0_aadd_2_a76.extended_lut = "off";
defparam fp_functions_0_aadd_2_a76.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a81(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a81_sumout),
	.cout(fp_functions_0_aadd_2_a82),
	.shareout());
defparam fp_functions_0_aadd_2_a81.extended_lut = "off";
defparam fp_functions_0_aadd_2_a81.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a86(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a86_sumout),
	.cout(fp_functions_0_aadd_2_a87),
	.shareout());
defparam fp_functions_0_aadd_2_a86.extended_lut = "off";
defparam fp_functions_0_aadd_2_a86.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a91(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a91_sumout),
	.cout(fp_functions_0_aadd_2_a92),
	.shareout());
defparam fp_functions_0_aadd_2_a91.extended_lut = "off";
defparam fp_functions_0_aadd_2_a91.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a96(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a96_sumout),
	.cout(fp_functions_0_aadd_2_a97),
	.shareout());
defparam fp_functions_0_aadd_2_a96.extended_lut = "off";
defparam fp_functions_0_aadd_2_a96.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_2_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a101(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a101_sumout),
	.cout(fp_functions_0_aadd_2_a102),
	.shareout());
defparam fp_functions_0_aadd_2_a101.extended_lut = "off";
defparam fp_functions_0_aadd_2_a101.lut_mask = 64'h0000000011116666;
defparam fp_functions_0_aadd_2_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a106(
	.dataa(!fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(!fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a106_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a106.extended_lut = "off";
defparam fp_functions_0_aadd_2_a106.lut_mask = 64'h0000000000006666;
defparam fp_functions_0_aadd_2_a106.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_5_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a6_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a5_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC0_uid62_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC0_uid62_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid62_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "00000000000000000000000000000000BFCB5221CD1082360385F58AAEDB6598";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a6_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_8_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_10_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[24]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a1_sumout),
	.cout(fp_functions_0_aadd_10_a2),
	.shareout());
defparam fp_functions_0_aadd_10_a1.extended_lut = "off";
defparam fp_functions_0_aadd_10_a1.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a6_sumout),
	.cout(fp_functions_0_aadd_10_a7),
	.shareout());
defparam fp_functions_0_aadd_10_a6.extended_lut = "off";
defparam fp_functions_0_aadd_10_a6.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[26]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a11_sumout),
	.cout(fp_functions_0_aadd_10_a12),
	.shareout());
defparam fp_functions_0_aadd_10_a11.extended_lut = "off";
defparam fp_functions_0_aadd_10_a11.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[27]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a16_sumout),
	.cout(fp_functions_0_aadd_10_a17),
	.shareout());
defparam fp_functions_0_aadd_10_a16.extended_lut = "off";
defparam fp_functions_0_aadd_10_a16.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[28]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a21_sumout),
	.cout(fp_functions_0_aadd_10_a22),
	.shareout());
defparam fp_functions_0_aadd_10_a21.extended_lut = "off";
defparam fp_functions_0_aadd_10_a21.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[29]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a26_sumout),
	.cout(fp_functions_0_aadd_10_a27),
	.shareout());
defparam fp_functions_0_aadd_10_a26.extended_lut = "off";
defparam fp_functions_0_aadd_10_a26.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a31_sumout),
	.cout(fp_functions_0_aadd_10_a32),
	.shareout());
defparam fp_functions_0_aadd_10_a31.extended_lut = "off";
defparam fp_functions_0_aadd_10_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_10_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_10_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_10_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_10_a36_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_10_a36.extended_lut = "off";
defparam fp_functions_0_aadd_10_a36.lut_mask = 64'h0000000000000000;
defparam fp_functions_0_aadd_10_a36.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout,fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout,
fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.ax_width = 12;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.ay_scan_in_width = 12;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.operation_mode = "m18x18_full";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.result_a_width = 24;
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.signed_max = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "0000000000000000000000000000000061E846A22F6F92639284430B2579B586";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "E16E0AA904653A99F52E85CFD4E0ECBDA58330823E9F8B8D601C8C81DD2FC839";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "E283D1FC00DB63CC28D4F74562ECAC36A43DC0219DE86D49EBD8E6835D88264D";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "E8E54C733023FD8C5E4726A6F3C3B0C7D4E24904E73E681780837088975DE957";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "B6E887B4B76E38D7590B0B2E43E24BF8F1142F42E8BBCA22440E36BE7FF783D1";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "94E502CD326410624F7B44A6A06F94CCA60D4F2B1AC689417D0419C4222244BD";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "8DB601A9CEC80A8110D3287641645D2DC7FCDA4C0654F72A7CA80AFD41417D09";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "8392AACE01DAACFF35631AB9D59D634CF803C6DAAB6700E6D6CFF9A980D58351";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "807199A5556CCF00F329ACC033567F2655556B6CCC78001E325AAD31FFCCAA61";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "800F879CCCDA5AAAA5B230FFF0CD2A4899998C70F07FFFFE0E399B6B55693381";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "2AAAD529696C933339C3C0FFF03CE6DA4B4B5AD5AAD55554AB52D24D998E3C01";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "66664C9B24DA49696B56AA555AA94B6CC738C63399CCCCCD99364924B4A56AAB";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "1E1E3C78E3C638E718CE66333664D9253F07C1F0783C3C3C78F1C71C739CE667";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "01FE03F81FC1F81F07C1E1F0F1E3C71CFF003FF007FC03FC07F03F03F07C1E1F";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "0001FFF8003FF800FFC01FF00FE03F0300FFFFF00003FFFC000FFF000FFC01FF";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "00000007FFFFF800003FFFF0001FFF00FFFFFFF000000003FFFFFF000003FFFF";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "00000000000007FFFFFFFFF0000000FFFFFFFFF000000000000000FFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "00000000000000000000000FFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC1_uid65_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fp_functions_0|memoryC1_uid65_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid65_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai768_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.address_width = 3;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.data_width = 1;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_address = 0;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_bit_number = 15;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.init_file = "none";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.last_address = 4;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_depth = 5;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_name = "fp_functions_0|redist7_yforpe_uid36_fpsqrttest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama15";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_width = 16;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1121_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1121_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1121_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a7_a_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_10_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!a[23]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_10_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_10_a42.extended_lut = "off";
defparam fp_functions_0_aadd_10_a42.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_10_a42.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_3_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_6_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a8_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a0_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a1_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a2_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a3_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a4_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a5_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a6_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a7_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a8_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a9_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a10_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a11_a_aq));
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai780_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai780_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai780_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a0_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a1_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a2_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a3_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a3_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai481_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist8_yaddr_uid35_fpsqrttest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a9_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "0000000000000000000000000000000001CEDD9304F7515E90834CC4CCEFE2F6";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "AC44C29DF2D1C8BC08CCBAFF4BB7B9C74E5D7A31458A8CC01F04C60A906635DB";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "3FF12EE758C74FD278FB1D98460289408B9E2D25912B55754AD21D46AFD93925";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "47798C899C1A6D24AD52AA35249187C00C1071C619CC66666C9B696BD5556B6C";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "787E0F0E1F1C71C7319CCCD9B6DAD56AF01F81F81E0F87878F1C718CE6664DB6";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "7F800FF01FE07E07C1E0F0E1C71CE673001FFE001FF007F80FE07E0F07878E38";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "7FFFF0001FFF8007FE00FF01F81F0783001FFFFFE00007FFF0007FF007F80FC0";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "7FFFFFFFE0000007FFFF0001FFE007FCFFE00000000007FFFFFF800007FFF000";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "7FFFFFFFFFFFFFF800000001FFFFF80000000000000007FFFFFFFFFFF8000000";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "800000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFE00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a_a23_a_a_wirecell_combout,a[22],a[21],a[20],a[19],a[18],a[17],a[16]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Sqrt_altera_fp_functions_191_wi5kdgi_memoryC2_uid68_sqrtTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC2_uid68_sqrtTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid68_sqrtTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a4_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a5_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a6_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a7_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a8_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a9_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a10_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a11_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a12_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a13_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a14_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a15_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_4_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a0_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a1_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a2_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a3_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_1_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_1_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a10_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a4_a(
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a4_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a5_a(
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a5_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a6_a(
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a6_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a7_a(
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a7_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a8_a(
	.clk(clk),
	.d(a[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a8_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a9_a(
	.clk(clk),
	.d(a[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a9_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a10_a(
	.clk(clk),
	.d(a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a10_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a11_a(
	.clk(clk),
	.d(a[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a11_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a12_a(
	.clk(clk),
	.d(a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a12_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a13_a(
	.clk(clk),
	.d(a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a13_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a14_a(
	.clk(clk),
	.d(a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a14_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a15_a(
	.clk(clk),
	.d(a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a15_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a0_a(
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a0_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a1_a(
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a1_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a2_a(
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a2_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a3_a(
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a3_a_aq));
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_delay_0_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai493_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai493_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai493_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a11_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_2_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a12_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a13_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_afracSel_uid48_fpSqrtTest_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a1_a_aq));
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a14_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_anegZero_uid59_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracSel_uid48_fpSqrtTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aMux_1_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_afracSel_uid48_fpSqrtTest_q_a1_a_aq));
defparam fp_functions_0_afracSel_uid48_fpSqrtTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_afracSel_uid48_fpSqrtTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anegZero_uid59_fpSqrtTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anegZero_uid59_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_anegZero_uid59_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_anegZero_uid59_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_9_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracXIsZero_uid15_fpSqrtTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_10_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid15_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid15_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid15_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a(
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_0_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aMux_32_a2(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_32_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_32_a2.extended_lut = "off";
defparam fp_functions_0_aMux_32_a2.lut_mask = 64'h1515151515151515;
defparam fp_functions_0_aMux_32_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_31_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_31_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_31_a0.extended_lut = "off";
defparam fp_functions_0_aMux_31_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_31_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_30_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_30_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_30_a0.extended_lut = "off";
defparam fp_functions_0_aMux_30_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_30_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_29_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_29_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_29_a0.extended_lut = "off";
defparam fp_functions_0_aMux_29_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_29_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_28_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_28_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_28_a0.extended_lut = "off";
defparam fp_functions_0_aMux_28_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_28_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_27_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_27_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_27_a0.extended_lut = "off";
defparam fp_functions_0_aMux_27_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_27_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_26_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_26_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_26_a0.extended_lut = "off";
defparam fp_functions_0_aMux_26_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_26_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_25_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_25_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_25_a0.extended_lut = "off";
defparam fp_functions_0_aMux_25_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_25_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_24_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_24_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_24_a0.extended_lut = "off";
defparam fp_functions_0_aMux_24_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_24_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_23_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_23_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_23_a0.extended_lut = "off";
defparam fp_functions_0_aMux_23_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_23_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_22_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_22_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_22_a0.extended_lut = "off";
defparam fp_functions_0_aMux_22_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_22_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_21_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_21_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_21_a0.extended_lut = "off";
defparam fp_functions_0_aMux_21_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_21_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_20_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_20_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_20_a0.extended_lut = "off";
defparam fp_functions_0_aMux_20_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_20_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_19_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_19_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_19_a0.extended_lut = "off";
defparam fp_functions_0_aMux_19_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_19_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_18_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_18_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_18_a0.extended_lut = "off";
defparam fp_functions_0_aMux_18_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_18_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_17_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_17_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_17_a0.extended_lut = "off";
defparam fp_functions_0_aMux_17_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_17_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_16_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_16_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_16_a0.extended_lut = "off";
defparam fp_functions_0_aMux_16_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_16_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_15_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_15_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_15_a0.extended_lut = "off";
defparam fp_functions_0_aMux_15_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_15_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_14_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_14_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_14_a0.extended_lut = "off";
defparam fp_functions_0_aMux_14_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_14_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_13_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_13_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_13_a0.extended_lut = "off";
defparam fp_functions_0_aMux_13_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_13_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_12_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_12_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_12_a0.extended_lut = "off";
defparam fp_functions_0_aMux_12_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_12_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_11_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_11_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_11_a0.extended_lut = "off";
defparam fp_functions_0_aMux_11_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_11_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_10_a0(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist5_fracRPostProcessings_uid39_fpSqrtTest_b_1_q_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_10_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_10_a0.extended_lut = "off";
defparam fp_functions_0_aMux_10_a0.lut_mask = 64'h0404040404040404;
defparam fp_functions_0_aMux_10_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a2(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a2.extended_lut = "off";
defparam fp_functions_0_aMux_9_a2.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a3(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a3.extended_lut = "off";
defparam fp_functions_0_aMux_9_a3.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a4(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a4.extended_lut = "off";
defparam fp_functions_0_aMux_9_a4.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a5(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a5.extended_lut = "off";
defparam fp_functions_0_aMux_9_a5.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a6(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a6.extended_lut = "off";
defparam fp_functions_0_aMux_9_a6.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a7(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a7.extended_lut = "off";
defparam fp_functions_0_aMux_9_a7.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a8(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a8.extended_lut = "off";
defparam fp_functions_0_aMux_9_a8.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a9(
	.dataa(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracSel_uid48_fpSqrtTest_q_16_adelay_signals_a0_a_a1_a_aq),
	.datac(!fp_functions_0_aredist3_expRR_uid51_fpSqrtTest_b_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a9.extended_lut = "off";
defparam fp_functions_0_aMux_9_a9.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_aMux_9_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a6_a_a0_a_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a36_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a37_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a38_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_lowRangeB_uid76_invPolyEval_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid78_invPolyEval_o_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ch_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1568_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1568_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai1568_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1410_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1410_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1410_a0.extended_lut = "off";
defparam fp_functions_0_ai1410_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai1410_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aexpRMux_uid31_fpSqrtTest_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1568_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1568_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1568_a0.extended_lut = "off";
defparam fp_functions_0_ai1568_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai1568_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1568_a1(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1568_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1568_a1.extended_lut = "off";
defparam fp_functions_0_ai1568_a1.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai1568_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1568_a2(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1568_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1568_a2.extended_lut = "off";
defparam fp_functions_0_ai1568_a2.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai1568_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_wraddr_q_a3_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11(
	.dataa(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a1_combout),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a0_combout),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a2_combout),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_cmp_b_a0_a_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11.lut_mask = 64'h0008000800080008;
defparam fp_functions_0_areduce_nor_11.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1140_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1109_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1109_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1109_a0.extended_lut = "off";
defparam fp_functions_0_ai1109_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai1109_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid90_pT2_uid81_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1424_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1424_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1424_a0.extended_lut = "off";
defparam fp_functions_0_ai1424_a0.lut_mask = 64'h6666666666666666;
defparam fp_functions_0_ai1424_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_8_a0(
	.dataa(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_8_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_8_a0.extended_lut = "off";
defparam fp_functions_0_aadd_8_a0.lut_mask = 64'h6969696969696969;
defparam fp_functions_0_aadd_8_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_8_a1(
	.dataa(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_8_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_8_a1.extended_lut = "off";
defparam fp_functions_0_aadd_8_a1.lut_mask = 64'h1E781E781E781E78;
defparam fp_functions_0_aadd_8_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_8_a2(
	.dataa(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a_aq),
	.datae(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_8_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_8_a2.extended_lut = "off";
defparam fp_functions_0_aadd_8_a2.lut_mask = 64'h01FE07F801FE07F8;
defparam fp_functions_0_aadd_8_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1140_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1140_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1140_a0.extended_lut = "off";
defparam fp_functions_0_ai1140_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai1140_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_5(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_5_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_5.extended_lut = "off";
defparam fp_functions_0_areduce_nor_5.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_8(
	.dataa(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist10_expRMux_uid31_fpSqrtTest_q_16_rdcnt_i_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_8_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_8.extended_lut = "off";
defparam fp_functions_0_areduce_nor_8.lut_mask = 64'h0008000800080008;
defparam fp_functions_0_areduce_nor_8.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_memoryC2_uid68_sqrtTables_lutmem_r_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid87_pT1_uid75_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai799_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai768_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai768_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai768_a0.extended_lut = "off";
defparam fp_functions_0_ai768_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai768_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_yForPe_uid36_fpSqrtTest_b_3_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq));
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1121_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1121_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1121_a0.extended_lut = "off";
defparam fp_functions_0_ai1121_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai1121_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1121_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1121_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1121_a1.extended_lut = "off";
defparam fp_functions_0_ai1121_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai1121_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1121_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1121_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1121_a2.extended_lut = "off";
defparam fp_functions_0_ai1121_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai1121_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai799_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai799_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai799_a0.extended_lut = "off";
defparam fp_functions_0_ai799_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai799_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_3(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_3_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_3.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6(
	.dataa(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist9_yAddr_uid35_fpSqrtTest_b_14_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai780_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai780_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai780_a0.extended_lut = "off";
defparam fp_functions_0_ai780_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai780_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai780_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai780_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai780_a1.extended_lut = "off";
defparam fp_functions_0_ai780_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai780_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai780_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai780_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai780_a2.extended_lut = "off";
defparam fp_functions_0_ai780_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai780_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai513_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(a[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai481_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai481_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai481_a0.extended_lut = "off";
defparam fp_functions_0_ai481_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai481_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(a[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(a[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4(
	.dataa(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist7_yForPe_uid36_fpSqrtTest_b_10_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai513_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai513_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai513_a0.extended_lut = "off";
defparam fp_functions_0_ai513_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai513_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai493_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai493_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai493_a0.extended_lut = "off";
defparam fp_functions_0_ai493_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai493_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai493_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai493_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai493_a1.extended_lut = "off";
defparam fp_functions_0_ai493_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai493_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai493_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai493_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai493_a2.extended_lut = "off";
defparam fp_functions_0_ai493_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai493_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_2(
	.dataa(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_2_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_2.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_2.shared_arith = "off";

fourteennm_ff fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1741_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a_aq));
defparam fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aMux_1_a0(
	.dataa(!fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_afracXIsZero_uid15_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_1_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_1_a0.extended_lut = "off";
defparam fp_functions_0_aMux_1_a0.lut_mask = 64'h10FA10FA10FA10FA;
defparam fp_functions_0_aMux_1_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1741_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_afracSel_uid48_fpSqrtTest_q_a0_a_aq),
	.datad(!fp_functions_0_aMux_1_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1741_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1741_a0.extended_lut = "off";
defparam fp_functions_0_ai1741_a0.lut_mask = 64'h7F5D7F5D7F5D7F5D;
defparam fp_functions_0_ai1741_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_1_a1(
	.dataa(!fp_functions_0_aexpXIsMax_uid14_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_1_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_1_a1.extended_lut = "off";
defparam fp_functions_0_aMux_1_a1.lut_mask = 64'h7171717171717171;
defparam fp_functions_0_aMux_1_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a(
	.dataa(!fp_functions_0_aredist11_signX_uid7_fpSqrtTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcZ_x_uid13_fpSqrtTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_anegZero_uid59_fpSqrtTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_9_a0(
	.dataa(!a[24]),
	.datab(!a[23]),
	.datac(!a[25]),
	.datad(!a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_9_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_9_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_9_a0.lut_mask = 64'h0001000100010001;
defparam fp_functions_0_areduce_nor_9_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_9(
	.dataa(!a[27]),
	.datab(!a[28]),
	.datac(!a[29]),
	.datad(!a[30]),
	.datae(!fp_functions_0_areduce_nor_9_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_9_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_9.extended_lut = "off";
defparam fp_functions_0_areduce_nor_9.lut_mask = 64'h0000000100000001;
defparam fp_functions_0_areduce_nor_9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a0(
	.dataa(!a[4]),
	.datab(!a[0]),
	.datac(!a[1]),
	.datad(!a[2]),
	.datae(!a[3]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_10_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a1(
	.dataa(!a[6]),
	.datab(!a[7]),
	.datac(!a[8]),
	.datad(!a[9]),
	.datae(!a[10]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a1.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_10_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a2(
	.dataa(!a[18]),
	.datab(!a[19]),
	.datac(!a[20]),
	.datad(!a[21]),
	.datae(!a[22]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a2.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_10_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a3(
	.dataa(!a[16]),
	.datab(!a[17]),
	.datac(!a[12]),
	.datad(!a[13]),
	.datae(!a[14]),
	.dataf(!a[15]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a3.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_areduce_nor_10_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10(
	.dataa(!a[5]),
	.datab(!a[11]),
	.datac(!fp_functions_0_areduce_nor_10_a0_combout),
	.datad(!fp_functions_0_areduce_nor_10_a1_combout),
	.datae(!fp_functions_0_areduce_nor_10_a2_combout),
	.dataf(!fp_functions_0_areduce_nor_10_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10.lut_mask = 64'h0000000000000008;
defparam fp_functions_0_areduce_nor_10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a0(
	.dataa(!a[24]),
	.datab(!a[23]),
	.datac(!a[25]),
	.datad(!a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_0_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0(
	.dataa(!a[27]),
	.datab(!a[28]),
	.datac(!a[29]),
	.datad(!a[30]),
	.datae(!fp_functions_0_areduce_nor_0_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0.lut_mask = 64'h0000800000008000;
defparam fp_functions_0_areduce_nor_0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0(
	.dataa(!a[23]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fp_functions_0_aredist8_yAddr_uid35_fpSqrtTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_a0.shared_arith = "off";

fourteennm_lcell_comb a_a23_a_a_wirecell(
	.dataa(!a[23]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(a_a23_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam a_a23_a_a_wirecell.extended_lut = "off";
defparam a_a23_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam a_a23_a_a_wirecell.shared_arith = "off";

assign q[22] = fp_functions_0_aMux_10_a0_combout;

assign q[21] = fp_functions_0_aMux_11_a0_combout;

assign q[20] = fp_functions_0_aMux_12_a0_combout;

assign q[19] = fp_functions_0_aMux_13_a0_combout;

assign q[18] = fp_functions_0_aMux_14_a0_combout;

assign q[17] = fp_functions_0_aMux_15_a0_combout;

assign q[16] = fp_functions_0_aMux_16_a0_combout;

assign q[15] = fp_functions_0_aMux_17_a0_combout;

assign q[14] = fp_functions_0_aMux_18_a0_combout;

assign q[13] = fp_functions_0_aMux_19_a0_combout;

assign q[12] = fp_functions_0_aMux_20_a0_combout;

assign q[11] = fp_functions_0_aMux_21_a0_combout;

assign q[10] = fp_functions_0_aMux_22_a0_combout;

assign q[9] = fp_functions_0_aMux_23_a0_combout;

assign q[8] = fp_functions_0_aMux_24_a0_combout;

assign q[7] = fp_functions_0_aMux_25_a0_combout;

assign q[6] = fp_functions_0_aMux_26_a0_combout;

assign q[5] = fp_functions_0_aMux_27_a0_combout;

assign q[4] = fp_functions_0_aMux_28_a0_combout;

assign q[3] = fp_functions_0_aMux_29_a0_combout;

assign q[2] = fp_functions_0_aMux_30_a0_combout;

assign q[1] = fp_functions_0_aMux_31_a0_combout;

assign q[0] = fp_functions_0_aMux_32_a2_combout;

assign q[23] = fp_functions_0_aMux_9_a2_combout;

assign q[24] = fp_functions_0_aMux_9_a3_combout;

assign q[25] = fp_functions_0_aMux_9_a4_combout;

assign q[26] = fp_functions_0_aMux_9_a5_combout;

assign q[27] = fp_functions_0_aMux_9_a6_combout;

assign q[28] = fp_functions_0_aMux_9_a7_combout;

assign q[29] = fp_functions_0_aMux_9_a8_combout;

assign q[30] = fp_functions_0_aMux_9_a9_combout;

assign q[31] = fp_functions_0_aredist2_negZero_uid59_fpSqrtTest_q_16_adelay_signals_a0_a_a0_a_aq;

endmodule
