module ItoF (
	input clk,
    input areset,
    input en,
    input signed [31:0] a,
    output logic [31:0] q 
);

    logic [31:0] pip0, pip1, pip2, pip3, pip4;
    int in;
    shortreal out;

    assign q = en ? pip4 : '0;
    always_comb begin 
        in = a;
        out = shortreal'(in);
    end

    always_ff @( posedge clk, posedge rst ) begin : internal_pipe
        if (rst) begin
            pip0 <= '0;
            pip1 <= '0;
            pip2 <= '0;
            pip3 <= '0;
            pip4 <= '0;

        end else begin
            if (en) begin
                pip0 <= $shortrealtobits(out);
                pip1 <= pip0;
                pip2 <= pip1;
                pip3 <= pip2;
                pip4 <= pip3;
            end else begin
                pip0 <= '0;
                pip1 <= '0;
                pip2 <= '0;
                pip3 <= '0;
                pip4 <= '0;
            end
                
        end
        
    end
endmodule