// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/20/2021 21:13:45"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Fix_Mul (
	result,
	clk,
	en,
	rst,
	b,
	a)/* synthesis synthesis_greybox=0 */;
output 	[63:0] result;
input 	clk;
input 	[0:0] en;
input 	rst;
input 	[31:0] b;
input 	[31:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fxp_functions_0_aadd_0_a1_sumout;
wire fxp_functions_0_aadd_0_a2;
wire fxp_functions_0_aadd_0_a6_sumout;
wire fxp_functions_0_aadd_0_a7;
wire fxp_functions_0_aadd_0_a11_sumout;
wire fxp_functions_0_aadd_0_a12;
wire fxp_functions_0_aadd_0_a16_sumout;
wire fxp_functions_0_aadd_0_a17;
wire fxp_functions_0_aadd_0_a21_sumout;
wire fxp_functions_0_aadd_0_a22;
wire fxp_functions_0_aadd_0_a26_sumout;
wire fxp_functions_0_aadd_0_a27;
wire fxp_functions_0_aadd_0_a31_sumout;
wire fxp_functions_0_aadd_0_a32;
wire fxp_functions_0_aadd_0_a36_sumout;
wire fxp_functions_0_aadd_0_a37;
wire fxp_functions_0_aadd_0_a41_sumout;
wire fxp_functions_0_aadd_0_a42;
wire fxp_functions_0_aadd_0_a46_sumout;
wire fxp_functions_0_aadd_0_a47;
wire fxp_functions_0_aadd_0_a51_sumout;
wire fxp_functions_0_aadd_0_a52;
wire fxp_functions_0_aadd_0_a56_sumout;
wire fxp_functions_0_aadd_0_a57;
wire fxp_functions_0_aadd_0_a61_sumout;
wire fxp_functions_0_aadd_0_a62;
wire fxp_functions_0_aadd_0_a66_sumout;
wire fxp_functions_0_aadd_0_a67;
wire fxp_functions_0_aadd_0_a71_sumout;
wire fxp_functions_0_aadd_0_a72;
wire fxp_functions_0_aadd_0_a76_sumout;
wire fxp_functions_0_aadd_0_a77;
wire fxp_functions_0_aadd_0_a81_sumout;
wire fxp_functions_0_aadd_0_a82;
wire fxp_functions_0_aadd_0_a86_sumout;
wire fxp_functions_0_aadd_0_a87;
wire fxp_functions_0_aadd_0_a91_sumout;
wire fxp_functions_0_aadd_0_a92;
wire fxp_functions_0_aadd_0_a96_sumout;
wire fxp_functions_0_aadd_0_a97;
wire fxp_functions_0_aadd_0_a101_sumout;
wire fxp_functions_0_aadd_0_a102;
wire fxp_functions_0_aadd_0_a106_sumout;
wire fxp_functions_0_aadd_0_a107;
wire fxp_functions_0_aadd_0_a111_sumout;
wire fxp_functions_0_aadd_0_a112;
wire fxp_functions_0_aadd_0_a116_sumout;
wire fxp_functions_0_aadd_0_a117;
wire fxp_functions_0_aadd_0_a121_sumout;
wire fxp_functions_0_aadd_0_a122;
wire fxp_functions_0_aadd_0_a126_sumout;
wire fxp_functions_0_aadd_0_a127;
wire fxp_functions_0_aadd_0_a131_sumout;
wire fxp_functions_0_aadd_0_a132;
wire fxp_functions_0_aadd_0_a136_sumout;
wire fxp_functions_0_aadd_0_a137;
wire fxp_functions_0_aadd_0_a141_sumout;
wire fxp_functions_0_aadd_0_a142;
wire fxp_functions_0_aadd_0_a146_sumout;
wire fxp_functions_0_aadd_0_a147;
wire fxp_functions_0_aadd_0_a151_sumout;
wire fxp_functions_0_aadd_0_a152;
wire fxp_functions_0_aadd_0_a156_sumout;
wire fxp_functions_0_aadd_0_a157;
wire fxp_functions_0_aadd_0_a161_sumout;
wire fxp_functions_0_aadd_0_a162;
wire fxp_functions_0_aadd_0_a166_sumout;
wire fxp_functions_0_aadd_0_a167;
wire fxp_functions_0_aadd_0_a171_sumout;
wire fxp_functions_0_aadd_0_a172;
wire fxp_functions_0_aadd_0_a176_sumout;
wire fxp_functions_0_aadd_0_a177;
wire fxp_functions_0_aadd_0_a181_sumout;
wire fxp_functions_0_aadd_0_a182;
wire fxp_functions_0_aadd_0_a186_sumout;
wire fxp_functions_0_aadd_0_a187;
wire fxp_functions_0_aadd_0_a191_sumout;
wire fxp_functions_0_aadd_0_a192;
wire fxp_functions_0_aadd_0_a196_sumout;
wire fxp_functions_0_aadd_0_a197;
wire fxp_functions_0_aadd_0_a201_sumout;
wire fxp_functions_0_aadd_0_a202;
wire fxp_functions_0_aadd_0_a206_sumout;
wire fxp_functions_0_aadd_0_a207;
wire fxp_functions_0_aadd_0_a211_sumout;
wire fxp_functions_0_aadd_0_a212;
wire fxp_functions_0_aadd_0_a216_sumout;
wire fxp_functions_0_aadd_0_a217;
wire fxp_functions_0_aadd_0_a221_sumout;
wire fxp_functions_0_aadd_0_a222;
wire fxp_functions_0_aadd_0_a226_sumout;
wire fxp_functions_0_amultiplier_im8_cma_s0_a0_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a1_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a2_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a3_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a4_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a5_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a6_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a7_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a8_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a9_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a10_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a11_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a12_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a13_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a14_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a15_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a16_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a17_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a18_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a19_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a20_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a21_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a22_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a23_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a24_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a25_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a26_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a27_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a28_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a29_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a30_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a31_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a32_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a33_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a34_a;
wire fxp_functions_0_amultiplier_im8_cma_s0_a35_a;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a0_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a1_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a2_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a3_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a4_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a5_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a6_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a7_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a8_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a9_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a10_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a11_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a12_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a13_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a14_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a15_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a16_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a17_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a18_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a19_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a20_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a21_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a22_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a23_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a24_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a25_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a26_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a27_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a28_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a29_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a30_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a31_a;
wire fxp_functions_0_amultiplier_ma3_cma_s0_a32_a;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA33;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA34;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA35;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_amultiplier_im0_cma_s0_a0_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a1_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a2_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a3_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a4_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a5_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a6_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a7_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a8_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a9_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a10_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a11_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a12_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a13_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a14_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a15_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a16_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a17_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a18_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a19_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a20_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a21_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a22_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a23_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a24_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a25_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a26_a;
wire fxp_functions_0_amultiplier_im0_cma_s0_a27_a;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA28;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA29;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA30;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA31;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA32;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA33;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA34;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA35;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a15_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a16_a_aq;
wire fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a17_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ena1_acombout;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a0_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a1_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a2_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a3_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a4_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a5_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a6_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a7_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a8_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a9_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a10_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a11_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a12_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a13_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a14_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a15_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a16_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a17_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a0_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a1_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a2_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a3_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a4_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a5_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a6_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a7_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a8_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a9_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a10_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a11_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a12_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a13_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a13_a_aq;

wire [63:0] fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus;
wire [63:0] fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus;
wire [63:0] fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus;

assign fxp_functions_0_amultiplier_im8_cma_s0_a0_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_amultiplier_im8_cma_s0_a1_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_amultiplier_im8_cma_s0_a2_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_amultiplier_im8_cma_s0_a3_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_amultiplier_im8_cma_s0_a4_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_amultiplier_im8_cma_s0_a5_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_amultiplier_im8_cma_s0_a6_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_amultiplier_im8_cma_s0_a7_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_amultiplier_im8_cma_s0_a8_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_amultiplier_im8_cma_s0_a9_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_amultiplier_im8_cma_s0_a10_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_amultiplier_im8_cma_s0_a11_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_amultiplier_im8_cma_s0_a12_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_amultiplier_im8_cma_s0_a13_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_amultiplier_im8_cma_s0_a14_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_amultiplier_im8_cma_s0_a15_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_amultiplier_im8_cma_s0_a16_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_amultiplier_im8_cma_s0_a17_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_amultiplier_im8_cma_s0_a18_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_amultiplier_im8_cma_s0_a19_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_amultiplier_im8_cma_s0_a20_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_amultiplier_im8_cma_s0_a21_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_amultiplier_im8_cma_s0_a22_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_amultiplier_im8_cma_s0_a23_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_amultiplier_im8_cma_s0_a24_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_amultiplier_im8_cma_s0_a25_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_amultiplier_im8_cma_s0_a26_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_amultiplier_im8_cma_s0_a27_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_amultiplier_im8_cma_s0_a28_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_amultiplier_im8_cma_s0_a29_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_amultiplier_im8_cma_s0_a30_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_amultiplier_im8_cma_s0_a31_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_amultiplier_im8_cma_s0_a32_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_amultiplier_im8_cma_s0_a33_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_amultiplier_im8_cma_s0_a34_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_amultiplier_im8_cma_s0_a35_a = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA36 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA37 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA38 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA39 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA40 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA41 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA42 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA43 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA44 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA45 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA46 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA47 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA48 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA49 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA50 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA51 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA52 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA53 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA54 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA55 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA56 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA57 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA58 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA59 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA60 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA61 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA62 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_amultiplier_im8_cma_DSP0_aDATAOUTA63 = fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_amultiplier_ma3_cma_s0_a0_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a1_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a2_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a3_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a4_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a5_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a6_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a7_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a8_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a9_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a10_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a11_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a12_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a13_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a14_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a15_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a16_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a17_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a18_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a19_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a20_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a21_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a22_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a23_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a24_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a25_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a26_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a27_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a28_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a29_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a30_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a31_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_amultiplier_ma3_cma_s0_a32_a = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA33 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA34 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA35 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA36 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA37 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA38 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA39 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA40 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA41 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA42 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA43 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA44 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA45 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA46 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA47 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA48 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA49 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA50 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA51 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA52 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA53 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA54 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA55 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA56 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA57 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA58 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA59 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA60 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA61 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA62 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_amultiplier_ma3_cma_DSP0_aDATAOUTA63 = fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_amultiplier_im0_cma_s0_a0_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_amultiplier_im0_cma_s0_a1_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_amultiplier_im0_cma_s0_a2_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_amultiplier_im0_cma_s0_a3_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_amultiplier_im0_cma_s0_a4_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_amultiplier_im0_cma_s0_a5_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_amultiplier_im0_cma_s0_a6_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_amultiplier_im0_cma_s0_a7_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_amultiplier_im0_cma_s0_a8_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_amultiplier_im0_cma_s0_a9_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_amultiplier_im0_cma_s0_a10_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_amultiplier_im0_cma_s0_a11_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_amultiplier_im0_cma_s0_a12_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_amultiplier_im0_cma_s0_a13_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_amultiplier_im0_cma_s0_a14_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_amultiplier_im0_cma_s0_a15_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_amultiplier_im0_cma_s0_a16_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_amultiplier_im0_cma_s0_a17_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_amultiplier_im0_cma_s0_a18_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_amultiplier_im0_cma_s0_a19_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_amultiplier_im0_cma_s0_a20_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_amultiplier_im0_cma_s0_a21_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_amultiplier_im0_cma_s0_a22_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_amultiplier_im0_cma_s0_a23_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_amultiplier_im0_cma_s0_a24_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_amultiplier_im0_cma_s0_a25_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_amultiplier_im0_cma_s0_a26_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_amultiplier_im0_cma_s0_a27_a = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA28 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA29 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA30 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA31 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA32 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA33 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA34 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA35 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA36 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA37 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA38 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA39 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA40 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA41 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA42 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA43 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA44 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA45 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA46 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA47 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA48 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA49 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA50 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA51 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA52 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA53 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA54 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA55 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA56 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA57 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA58 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA59 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA60 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA61 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA62 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_amultiplier_im0_cma_DSP0_aDATAOUTA63 = fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus[63];

fourteennm_lcell_comb fxp_functions_0_aadd_0_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a1_sumout),
	.cout(fxp_functions_0_aadd_0_a2),
	.shareout());
defparam fxp_functions_0_aadd_0_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a1.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a6_sumout),
	.cout(fxp_functions_0_aadd_0_a7),
	.shareout());
defparam fxp_functions_0_aadd_0_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a6.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a11_sumout),
	.cout(fxp_functions_0_aadd_0_a12),
	.shareout());
defparam fxp_functions_0_aadd_0_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a11.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a16_sumout),
	.cout(fxp_functions_0_aadd_0_a17),
	.shareout());
defparam fxp_functions_0_aadd_0_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a16.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a21_sumout),
	.cout(fxp_functions_0_aadd_0_a22),
	.shareout());
defparam fxp_functions_0_aadd_0_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a21.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a26_sumout),
	.cout(fxp_functions_0_aadd_0_a27),
	.shareout());
defparam fxp_functions_0_aadd_0_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a26.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a31_sumout),
	.cout(fxp_functions_0_aadd_0_a32),
	.shareout());
defparam fxp_functions_0_aadd_0_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a31.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a36_sumout),
	.cout(fxp_functions_0_aadd_0_a37),
	.shareout());
defparam fxp_functions_0_aadd_0_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a36.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a41_sumout),
	.cout(fxp_functions_0_aadd_0_a42),
	.shareout());
defparam fxp_functions_0_aadd_0_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a41.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a46_sumout),
	.cout(fxp_functions_0_aadd_0_a47),
	.shareout());
defparam fxp_functions_0_aadd_0_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a46.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a51_sumout),
	.cout(fxp_functions_0_aadd_0_a52),
	.shareout());
defparam fxp_functions_0_aadd_0_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a51.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a56_sumout),
	.cout(fxp_functions_0_aadd_0_a57),
	.shareout());
defparam fxp_functions_0_aadd_0_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a56.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a61_sumout),
	.cout(fxp_functions_0_aadd_0_a62),
	.shareout());
defparam fxp_functions_0_aadd_0_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a61.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a66_sumout),
	.cout(fxp_functions_0_aadd_0_a67),
	.shareout());
defparam fxp_functions_0_aadd_0_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a66.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a71_sumout),
	.cout(fxp_functions_0_aadd_0_a72),
	.shareout());
defparam fxp_functions_0_aadd_0_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a71.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a76_sumout),
	.cout(fxp_functions_0_aadd_0_a77),
	.shareout());
defparam fxp_functions_0_aadd_0_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a76.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a81_sumout),
	.cout(fxp_functions_0_aadd_0_a82),
	.shareout());
defparam fxp_functions_0_aadd_0_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a81.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a86_sumout),
	.cout(fxp_functions_0_aadd_0_a87),
	.shareout());
defparam fxp_functions_0_aadd_0_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a86.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a91_sumout),
	.cout(fxp_functions_0_aadd_0_a92),
	.shareout());
defparam fxp_functions_0_aadd_0_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a91.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a1_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a96_sumout),
	.cout(fxp_functions_0_aadd_0_a97),
	.shareout());
defparam fxp_functions_0_aadd_0_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a96.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a2_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a101_sumout),
	.cout(fxp_functions_0_aadd_0_a102),
	.shareout());
defparam fxp_functions_0_aadd_0_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a101.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a3_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a106_sumout),
	.cout(fxp_functions_0_aadd_0_a107),
	.shareout());
defparam fxp_functions_0_aadd_0_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a106.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a4_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a111_sumout),
	.cout(fxp_functions_0_aadd_0_a112),
	.shareout());
defparam fxp_functions_0_aadd_0_a111.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a111.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a111.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a5_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a116_sumout),
	.cout(fxp_functions_0_aadd_0_a117),
	.shareout());
defparam fxp_functions_0_aadd_0_a116.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a116.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a116.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a6_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a121_sumout),
	.cout(fxp_functions_0_aadd_0_a122),
	.shareout());
defparam fxp_functions_0_aadd_0_a121.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a121.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a121.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a7_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a126_sumout),
	.cout(fxp_functions_0_aadd_0_a127),
	.shareout());
defparam fxp_functions_0_aadd_0_a126.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a126.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a126.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a8_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a131_sumout),
	.cout(fxp_functions_0_aadd_0_a132),
	.shareout());
defparam fxp_functions_0_aadd_0_a131.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a131.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a131.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a9_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a136_sumout),
	.cout(fxp_functions_0_aadd_0_a137),
	.shareout());
defparam fxp_functions_0_aadd_0_a136.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a136.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a136.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a10_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a141_sumout),
	.cout(fxp_functions_0_aadd_0_a142),
	.shareout());
defparam fxp_functions_0_aadd_0_a141.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a141.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a141.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a146_sumout),
	.cout(fxp_functions_0_aadd_0_a147),
	.shareout());
defparam fxp_functions_0_aadd_0_a146.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a146.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a146.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a151_sumout),
	.cout(fxp_functions_0_aadd_0_a152),
	.shareout());
defparam fxp_functions_0_aadd_0_a151.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a151.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a151.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a156(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datad(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a156_sumout),
	.cout(fxp_functions_0_aadd_0_a157),
	.shareout());
defparam fxp_functions_0_aadd_0_a156.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a156.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_0_a156.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a161(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a157),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a161_sumout),
	.cout(fxp_functions_0_aadd_0_a162),
	.shareout());
defparam fxp_functions_0_aadd_0_a161.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a161.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a161.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a166(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a162),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a166_sumout),
	.cout(fxp_functions_0_aadd_0_a167),
	.shareout());
defparam fxp_functions_0_aadd_0_a166.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a166.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a166.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a171(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a167),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a171_sumout),
	.cout(fxp_functions_0_aadd_0_a172),
	.shareout());
defparam fxp_functions_0_aadd_0_a171.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a171.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a171.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a176(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a172),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a176_sumout),
	.cout(fxp_functions_0_aadd_0_a177),
	.shareout());
defparam fxp_functions_0_aadd_0_a176.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a176.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a176.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a181(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a177),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a181_sumout),
	.cout(fxp_functions_0_aadd_0_a182),
	.shareout());
defparam fxp_functions_0_aadd_0_a181.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a181.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a181.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a186(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a182),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a186_sumout),
	.cout(fxp_functions_0_aadd_0_a187),
	.shareout());
defparam fxp_functions_0_aadd_0_a186.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a186.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a186.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a191(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a187),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a191_sumout),
	.cout(fxp_functions_0_aadd_0_a192),
	.shareout());
defparam fxp_functions_0_aadd_0_a191.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a191.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a191.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a196(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a192),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a196_sumout),
	.cout(fxp_functions_0_aadd_0_a197),
	.shareout());
defparam fxp_functions_0_aadd_0_a196.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a196.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a196.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a201(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a197),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a201_sumout),
	.cout(fxp_functions_0_aadd_0_a202),
	.shareout());
defparam fxp_functions_0_aadd_0_a201.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a201.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a201.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a206(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a202),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a206_sumout),
	.cout(fxp_functions_0_aadd_0_a207),
	.shareout());
defparam fxp_functions_0_aadd_0_a206.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a206.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a206.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a211(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a207),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a211_sumout),
	.cout(fxp_functions_0_aadd_0_a212),
	.shareout());
defparam fxp_functions_0_aadd_0_a211.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a211.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a211.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a216(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a212),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a216_sumout),
	.cout(fxp_functions_0_aadd_0_a217),
	.shareout());
defparam fxp_functions_0_aadd_0_a216.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a216.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a216.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a221(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a217),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a221_sumout),
	.cout(fxp_functions_0_aadd_0_a222),
	.shareout());
defparam fxp_functions_0_aadd_0_a221.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a221.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_0_a221.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a226(
	.dataa(!fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_0_a222),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_0_a226_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_0_a226.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a226.lut_mask = 64'h0000000000005A5A;
defparam fxp_functions_0_aadd_0_a226.shared_arith = "off";

fourteennm_mac fxp_functions_0_amultiplier_im8_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a17_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a16_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a15_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a14_a_aq,
fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a13_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a12_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a11_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a10_a_aq,
fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a9_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a8_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a7_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a6_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a5_a_aq,
fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a4_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a3_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a2_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a1_a_aq,fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a17_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a16_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a15_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a14_a_aq,
fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a13_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a12_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a11_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a10_a_aq,
fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a9_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a8_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a7_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a6_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a5_a_aq,
fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a4_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a3_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a2_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a1_a_aq,fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_amultiplier_ma3_cma_ena1_acombout,fxp_functions_0_amultiplier_ma3_cma_ena1_acombout,fxp_functions_0_amultiplier_ma3_cma_ena1_acombout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_amultiplier_im8_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.ax_width = 18;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.ay_scan_in_width = 18;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.operation_mode = "m18x18_full";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.result_a_width = 36;
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.signed_max = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.signed_may = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_amultiplier_im8_cma_DSP0.use_chainadder = "false";

fourteennm_mac fxp_functions_0_amultiplier_ma3_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a17_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a16_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a15_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a14_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a13_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a12_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a11_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a10_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a9_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a8_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a7_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a6_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a5_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a4_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a3_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a2_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a1_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a13_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a12_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a11_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a10_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a9_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a8_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a7_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a6_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a5_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a4_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a3_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a2_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a1_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx({fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a17_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a16_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a15_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a14_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a13_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a12_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a11_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a10_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a9_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a8_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a7_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a6_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a5_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a4_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a3_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a2_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a1_a_aq,fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a0_a_aq}),
	.by({gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a13_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a12_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a11_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a10_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a9_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a8_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a7_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a6_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a5_a_aq,
fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a4_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a3_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a2_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a1_a_aq,fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a0_a_aq}),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_amultiplier_ma3_cma_ena1_acombout,fxp_functions_0_amultiplier_ma3_cma_ena1_acombout,fxp_functions_0_amultiplier_ma3_cma_ena1_acombout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_amultiplier_ma3_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.ax_width = 18;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.ay_scan_in_width = 14;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.bx_clock = "0";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.bx_width = 18;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.by_clock = "0";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.by_width = 14;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.operation_mode = "m18x18_sumof2";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.result_a_width = 33;
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.signed_max = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.signed_may = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.signed_mby = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_amultiplier_ma3_cma_DSP0.use_chainadder = "false";

fourteennm_mac fxp_functions_0_amultiplier_im0_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a13_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a12_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a11_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a10_a_aq,
fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a9_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a8_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a7_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a6_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a5_a_aq,
fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a4_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a3_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a2_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a1_a_aq,fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a13_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a12_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a11_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a10_a_aq,
fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a9_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a8_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a7_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a6_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a5_a_aq,
fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a4_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a3_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a2_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a1_a_aq,fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_amultiplier_ma3_cma_ena1_acombout,fxp_functions_0_amultiplier_ma3_cma_ena1_acombout,fxp_functions_0_amultiplier_ma3_cma_ena1_acombout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_amultiplier_im0_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.ax_width = 14;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.ay_scan_in_width = 14;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.operation_mode = "m18x18_full";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.result_a_width = 28;
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.signed_max = "true";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.signed_may = "true";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_amultiplier_im0_cma_DSP0.use_chainadder = "false";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im8_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_ma3_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_amultiplier_im0_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(b[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(b[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(b[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(b[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(b[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(b[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(b[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(b[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(b[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(a[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(a[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(a[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a16_a(
	.clk(clk),
	.d(a[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a17_a(
	.clk(clk),
	.d(a[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im8_cma_ah_a0_a_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_amultiplier_ma3_cma_ena1(
	.dataa(!en[0]),
	.datab(!rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultiplier_ma3_cma_ena1_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultiplier_ma3_cma_ena1.extended_lut = "off";
defparam fxp_functions_0_amultiplier_ma3_cma_ena1.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_amultiplier_ma3_cma_ena1.shared_arith = "off";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a0_a(
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a1_a(
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a2_a(
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a3_a(
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a4_a(
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a5_a(
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a6_a(
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a7_a(
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a8_a(
	.clk(clk),
	.d(a[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a9_a(
	.clk(clk),
	.d(a[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a10_a(
	.clk(clk),
	.d(a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a11_a(
	.clk(clk),
	.d(a[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a12_a(
	.clk(clk),
	.d(a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a13_a(
	.clk(clk),
	.d(a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a14_a(
	.clk(clk),
	.d(a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a15_a(
	.clk(clk),
	.d(a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a16_a(
	.clk(clk),
	.d(a[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a17_a(
	.clk(clk),
	.d(a[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a1_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a0_a(
	.clk(clk),
	.d(b[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a1_a(
	.clk(clk),
	.d(b[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a2_a(
	.clk(clk),
	.d(b[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a3_a(
	.clk(clk),
	.d(b[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a4_a(
	.clk(clk),
	.d(b[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a5_a(
	.clk(clk),
	.d(b[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a6_a(
	.clk(clk),
	.d(b[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a7_a(
	.clk(clk),
	.d(b[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a8_a(
	.clk(clk),
	.d(b[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a9_a(
	.clk(clk),
	.d(b[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a10_a(
	.clk(clk),
	.d(b[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a11_a(
	.clk(clk),
	.d(b[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a12_a(
	.clk(clk),
	.d(b[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a13_a(
	.clk(clk),
	.d(b[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a1_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(b[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(b[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(b[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(b[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(b[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(b[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(b[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(b[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(b[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(a[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(a[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(a[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(a[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(a[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(a[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(a[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(a[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(a[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_ma3_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(b[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(b[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(b[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(b[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(b[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(b[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(b[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(b[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(b[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(b[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(b[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(b[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(b[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(b[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(a[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(a[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(a[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(a[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(a[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(a[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(a[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(a[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(a[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultiplier_im0_cma_ah_a0_a_a13_a.power_up = "dont_care";

assign result[38] = fxp_functions_0_aadd_0_a101_sumout;

assign result[39] = fxp_functions_0_aadd_0_a106_sumout;

assign result[40] = fxp_functions_0_aadd_0_a111_sumout;

assign result[41] = fxp_functions_0_aadd_0_a116_sumout;

assign result[20] = fxp_functions_0_aadd_0_a11_sumout;

assign result[42] = fxp_functions_0_aadd_0_a121_sumout;

assign result[43] = fxp_functions_0_aadd_0_a126_sumout;

assign result[44] = fxp_functions_0_aadd_0_a131_sumout;

assign result[45] = fxp_functions_0_aadd_0_a136_sumout;

assign result[46] = fxp_functions_0_aadd_0_a141_sumout;

assign result[47] = fxp_functions_0_aadd_0_a146_sumout;

assign result[48] = fxp_functions_0_aadd_0_a151_sumout;

assign result[49] = fxp_functions_0_aadd_0_a156_sumout;

assign result[50] = fxp_functions_0_aadd_0_a161_sumout;

assign result[51] = fxp_functions_0_aadd_0_a166_sumout;

assign result[21] = fxp_functions_0_aadd_0_a16_sumout;

assign result[52] = fxp_functions_0_aadd_0_a171_sumout;

assign result[53] = fxp_functions_0_aadd_0_a176_sumout;

assign result[54] = fxp_functions_0_aadd_0_a181_sumout;

assign result[55] = fxp_functions_0_aadd_0_a186_sumout;

assign result[56] = fxp_functions_0_aadd_0_a191_sumout;

assign result[57] = fxp_functions_0_aadd_0_a196_sumout;

assign result[18] = fxp_functions_0_aadd_0_a1_sumout;

assign result[58] = fxp_functions_0_aadd_0_a201_sumout;

assign result[59] = fxp_functions_0_aadd_0_a206_sumout;

assign result[60] = fxp_functions_0_aadd_0_a211_sumout;

assign result[61] = fxp_functions_0_aadd_0_a216_sumout;

assign result[22] = fxp_functions_0_aadd_0_a21_sumout;

assign result[62] = fxp_functions_0_aadd_0_a221_sumout;

assign result[63] = fxp_functions_0_aadd_0_a226_sumout;

assign result[23] = fxp_functions_0_aadd_0_a26_sumout;

assign result[24] = fxp_functions_0_aadd_0_a31_sumout;

assign result[25] = fxp_functions_0_aadd_0_a36_sumout;

assign result[26] = fxp_functions_0_aadd_0_a41_sumout;

assign result[27] = fxp_functions_0_aadd_0_a46_sumout;

assign result[28] = fxp_functions_0_aadd_0_a51_sumout;

assign result[29] = fxp_functions_0_aadd_0_a56_sumout;

assign result[30] = fxp_functions_0_aadd_0_a61_sumout;

assign result[31] = fxp_functions_0_aadd_0_a66_sumout;

assign result[19] = fxp_functions_0_aadd_0_a6_sumout;

assign result[32] = fxp_functions_0_aadd_0_a71_sumout;

assign result[33] = fxp_functions_0_aadd_0_a76_sumout;

assign result[34] = fxp_functions_0_aadd_0_a81_sumout;

assign result[35] = fxp_functions_0_aadd_0_a86_sumout;

assign result[36] = fxp_functions_0_aadd_0_a91_sumout;

assign result[37] = fxp_functions_0_aadd_0_a96_sumout;

assign result[0] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a0_a_aq;

assign result[10] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a10_a_aq;

assign result[11] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a11_a_aq;

assign result[12] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a12_a_aq;

assign result[13] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a13_a_aq;

assign result[14] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a14_a_aq;

assign result[15] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a15_a_aq;

assign result[16] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a16_a_aq;

assign result[17] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a17_a_aq;

assign result[1] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a1_a_aq;

assign result[2] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a2_a_aq;

assign result[3] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a3_a_aq;

assign result[4] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a4_a_aq;

assign result[5] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a5_a_aq;

assign result[6] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a6_a_aq;

assign result[7] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a7_a_aq;

assign result[8] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a8_a_aq;

assign result[9] = fxp_functions_0_amultiplier_im8_cma_delay_adelay_signals_a0_a_a9_a_aq;

endmodule
