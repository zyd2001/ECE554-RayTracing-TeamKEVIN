module Float_Sub (
		input  wire        clk0,   //   clk0.clk
		input  wire        ena,    //    ena.ena
		input  wire        clr0,   //   clr0.reset
		input  wire        clr1,   //   clr1.reset
		output wire [31:0] result, // result.result
		input  wire [31:0] ax,     //     ax.ax
		input  wire [31:0] ay      //     ay.ay
	);
endmodule

