// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/20/2021 22:56:03"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Fix_Sqrt (
	result,
	clk,
	rst,
	en,
	radical)/* synthesis synthesis_greybox=0 */;
output 	[31:0] result;
input 	clk;
input 	rst;
input 	[0:0] en;
input 	[31:0] radical;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fxp_functions_0_aadd_32_a1_sumout;
wire fxp_functions_0_aadd_32_a2;
wire fxp_functions_0_aadd_32_a6_sumout;
wire fxp_functions_0_aadd_32_a7;
wire fxp_functions_0_aadd_32_a11_sumout;
wire fxp_functions_0_aadd_32_a12;
wire fxp_functions_0_aadd_32_a16_sumout;
wire fxp_functions_0_aadd_32_a17;
wire fxp_functions_0_aadd_32_a21_sumout;
wire fxp_functions_0_aadd_32_a22;
wire fxp_functions_0_aadd_32_a26_sumout;
wire fxp_functions_0_aadd_32_a27;
wire fxp_functions_0_aadd_32_a31_sumout;
wire fxp_functions_0_aadd_32_a32;
wire fxp_functions_0_aadd_32_a36_sumout;
wire fxp_functions_0_aadd_32_a37;
wire fxp_functions_0_aadd_32_a41_sumout;
wire fxp_functions_0_aadd_32_a42;
wire fxp_functions_0_aadd_32_a46_sumout;
wire fxp_functions_0_aadd_32_a47;
wire fxp_functions_0_aadd_32_a51_sumout;
wire fxp_functions_0_aadd_32_a52;
wire fxp_functions_0_aadd_32_a56_sumout;
wire fxp_functions_0_aadd_32_a57;
wire fxp_functions_0_aadd_32_a61_sumout;
wire fxp_functions_0_aadd_32_a62;
wire fxp_functions_0_aadd_32_a66_sumout;
wire fxp_functions_0_aadd_32_a67;
wire fxp_functions_0_aadd_32_a71_sumout;
wire fxp_functions_0_aadd_32_a72;
wire fxp_functions_0_aadd_32_a76_sumout;
wire fxp_functions_0_aadd_32_a77;
wire fxp_functions_0_aadd_32_a81_sumout;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aadd_31_a1_sumout;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a_aq;
wire fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a_aq;
wire fxp_functions_0_aadd_29_a1_sumout;
wire fxp_functions_0_aadd_31_a7_cout;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a_aq;
wire fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a_aq;
wire fxp_functions_0_aadd_29_a7_cout;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a18_a_aq;
wire fxp_functions_0_aadd_31_a12_cout;
wire fxp_functions_0_aadd_27_a1_sumout;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a_aq;
wire fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a_aq;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a17_a_aq;
wire fxp_functions_0_aadd_29_a12_cout;
wire fxp_functions_0_aadd_30_a1_sumout;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a17_a_aq;
wire fxp_functions_0_aadd_31_a17_cout;
wire fxp_functions_0_aadd_27_a7_cout;
wire fxp_functions_0_aadd_25_a1_sumout;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a_aq;
wire fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a_aq;
wire fxp_functions_0_aadd_28_a1_sumout;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a_aq;
wire fxp_functions_0_aadd_29_a17_cout;
wire fxp_functions_0_aadd_30_a6_sumout;
wire fxp_functions_0_aadd_30_a7;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a16_a_aq;
wire fxp_functions_0_aadd_31_a22_cout;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a16_a_aq;
wire fxp_functions_0_aadd_27_a12_cout;
wire fxp_functions_0_aadd_25_a7_cout;
wire fxp_functions_0_aadd_23_a1_sumout;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a_aq;
wire fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a_aq;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a_aq;
wire fxp_functions_0_aadd_28_a6_sumout;
wire fxp_functions_0_aadd_28_a7;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a_aq;
wire fxp_functions_0_aadd_29_a22_cout;
wire fxp_functions_0_aadd_30_a11_sumout;
wire fxp_functions_0_aadd_30_a12;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a15_a_aq;
wire fxp_functions_0_aadd_31_a27_cout;
wire fxp_functions_0_aadd_26_a1_sumout;
wire fxp_functions_0_aadd_27_a17_cout;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a15_a_aq;
wire fxp_functions_0_aadd_25_a12_cout;
wire fxp_functions_0_aadd_23_a7_cout;
wire fxp_functions_0_aadd_21_a1_sumout;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a_aq;
wire fxp_functions_0_aadd_26_a6_sumout;
wire fxp_functions_0_aadd_26_a7;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a_aq;
wire fxp_functions_0_aadd_28_a11_sumout;
wire fxp_functions_0_aadd_28_a12;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a_aq;
wire fxp_functions_0_aadd_29_a27_cout;
wire fxp_functions_0_aadd_30_a16_sumout;
wire fxp_functions_0_aadd_30_a17;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a14_a_aq;
wire fxp_functions_0_aadd_31_a32_cout;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a_aq;
wire fxp_functions_0_aadd_27_a22_cout;
wire fxp_functions_0_aadd_24_a1_sumout;
wire fxp_functions_0_aadd_25_a17_cout;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a14_a_aq;
wire fxp_functions_0_aadd_23_a12_cout;
wire fxp_functions_0_aadd_21_a7_cout;
wire fxp_functions_0_aadd_19_a1_sumout;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a_aq;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a_aq;
wire fxp_functions_0_aadd_26_a11_sumout;
wire fxp_functions_0_aadd_26_a12;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a_aq;
wire fxp_functions_0_aadd_28_a16_sumout;
wire fxp_functions_0_aadd_28_a17;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a_aq;
wire fxp_functions_0_aadd_29_a32_cout;
wire fxp_functions_0_aadd_30_a21_sumout;
wire fxp_functions_0_aadd_30_a22;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a13_a_aq;
wire fxp_functions_0_aadd_31_a37_cout;
wire fxp_functions_0_aadd_24_a6_sumout;
wire fxp_functions_0_aadd_24_a7;
wire fxp_functions_0_aadd_27_a27_cout;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a_aq;
wire fxp_functions_0_aadd_25_a22_cout;
wire fxp_functions_0_aadd_22_a1_sumout;
wire fxp_functions_0_aadd_23_a17_cout;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a13_a_aq;
wire fxp_functions_0_aadd_21_a12_cout;
wire fxp_functions_0_aadd_19_a7_cout;
wire fxp_functions_0_aadd_17_a1_sumout;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a_aq;
wire fxp_functions_0_aadd_24_a11_sumout;
wire fxp_functions_0_aadd_24_a12;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a_aq;
wire fxp_functions_0_aadd_26_a16_sumout;
wire fxp_functions_0_aadd_26_a17;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a_aq;
wire fxp_functions_0_aadd_28_a21_sumout;
wire fxp_functions_0_aadd_28_a22;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a_aq;
wire fxp_functions_0_aadd_29_a37_cout;
wire fxp_functions_0_aadd_30_a26_sumout;
wire fxp_functions_0_aadd_30_a27;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a12_a_aq;
wire fxp_functions_0_aadd_31_a42_cout;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a_aq;
wire fxp_functions_0_aadd_27_a32_cout;
wire fxp_functions_0_aadd_22_a6_sumout;
wire fxp_functions_0_aadd_22_a7;
wire fxp_functions_0_aadd_25_a27_cout;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a_aq;
wire fxp_functions_0_aadd_23_a22_cout;
wire fxp_functions_0_aadd_20_a1_sumout;
wire fxp_functions_0_aadd_21_a17_cout;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a12_a_aq;
wire fxp_functions_0_aadd_19_a12_cout;
wire fxp_functions_0_aadd_17_a7_cout;
wire fxp_functions_0_aadd_15_a1_sumout;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a_aq;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_24_a16_sumout;
wire fxp_functions_0_aadd_24_a17;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_26_a21_sumout;
wire fxp_functions_0_aadd_26_a22;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_28_a26_sumout;
wire fxp_functions_0_aadd_28_a27;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_29_a42_cout;
wire fxp_functions_0_aadd_30_a31_sumout;
wire fxp_functions_0_aadd_30_a32;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a11_a_aq;
wire fxp_functions_0_aadd_31_a47_cout;
wire fxp_functions_0_aadd_22_a11_sumout;
wire fxp_functions_0_aadd_22_a12;
wire fxp_functions_0_aadd_27_a37_cout;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_25_a32_cout;
wire fxp_functions_0_aadd_20_a6_sumout;
wire fxp_functions_0_aadd_20_a7;
wire fxp_functions_0_aadd_23_a27_cout;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_21_a22_cout;
wire fxp_functions_0_aadd_18_a1_sumout;
wire fxp_functions_0_aadd_19_a17_cout;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a11_a_aq;
wire fxp_functions_0_aadd_17_a12_cout;
wire fxp_functions_0_aadd_15_a7_cout;
wire fxp_functions_0_aadd_13_a1_sumout;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a_aq;
wire fxp_functions_0_aadd_22_a16_sumout;
wire fxp_functions_0_aadd_22_a17;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_24_a21_sumout;
wire fxp_functions_0_aadd_24_a22;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_26_a26_sumout;
wire fxp_functions_0_aadd_26_a27;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_28_a31_sumout;
wire fxp_functions_0_aadd_28_a32;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_29_a47_cout;
wire fxp_functions_0_aadd_30_a36_sumout;
wire fxp_functions_0_aadd_30_a37;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a10_a_aq;
wire fxp_functions_0_aadd_31_a52_cout;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_27_a42_cout;
wire fxp_functions_0_aadd_20_a11_sumout;
wire fxp_functions_0_aadd_20_a12;
wire fxp_functions_0_aadd_25_a37_cout;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_23_a32_cout;
wire fxp_functions_0_aadd_18_a6_sumout;
wire fxp_functions_0_aadd_18_a7;
wire fxp_functions_0_aadd_21_a27_cout;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_19_a22_cout;
wire fxp_functions_0_aadd_16_a1_sumout;
wire fxp_functions_0_aadd_17_a17_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a10_a_aq;
wire fxp_functions_0_aadd_15_a12_cout;
wire fxp_functions_0_aadd_13_a7_cout;
wire fxp_functions_0_aadd_11_a1_sumout;
wire fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_22_a21_sumout;
wire fxp_functions_0_aadd_22_a22;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_24_a26_sumout;
wire fxp_functions_0_aadd_24_a27;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_26_a31_sumout;
wire fxp_functions_0_aadd_26_a32;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_28_a36_sumout;
wire fxp_functions_0_aadd_28_a37;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_29_a52_cout;
wire fxp_functions_0_aadd_30_a41_sumout;
wire fxp_functions_0_aadd_30_a42;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a9_a_aq;
wire fxp_functions_0_aadd_31_a57_cout;
wire fxp_functions_0_aadd_20_a16_sumout;
wire fxp_functions_0_aadd_20_a17;
wire fxp_functions_0_aadd_27_a47_cout;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_25_a42_cout;
wire fxp_functions_0_aadd_18_a11_sumout;
wire fxp_functions_0_aadd_18_a12;
wire fxp_functions_0_aadd_23_a37_cout;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_21_a32_cout;
wire fxp_functions_0_aadd_16_a6_sumout;
wire fxp_functions_0_aadd_16_a7;
wire fxp_functions_0_aadd_19_a27_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_17_a22_cout;
wire fxp_functions_0_aadd_14_a1_sumout;
wire fxp_functions_0_aadd_15_a17_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a9_a_aq;
wire fxp_functions_0_aadd_13_a12_cout;
wire fxp_functions_0_aadd_11_a7_cout;
wire fxp_functions_0_aadd_9_a1_sumout;
wire fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a_aq;
wire fxp_functions_0_aadd_20_a21_sumout;
wire fxp_functions_0_aadd_20_a22;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_22_a26_sumout;
wire fxp_functions_0_aadd_22_a27;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_24_a31_sumout;
wire fxp_functions_0_aadd_24_a32;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_26_a36_sumout;
wire fxp_functions_0_aadd_26_a37;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_28_a41_sumout;
wire fxp_functions_0_aadd_28_a42;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_29_a57_cout;
wire fxp_functions_0_aadd_30_a46_sumout;
wire fxp_functions_0_aadd_30_a47;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a8_a_aq;
wire fxp_functions_0_aadd_31_a62_cout;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_27_a52_cout;
wire fxp_functions_0_aadd_18_a16_sumout;
wire fxp_functions_0_aadd_18_a17;
wire fxp_functions_0_aadd_25_a47_cout;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_23_a42_cout;
wire fxp_functions_0_aadd_16_a11_sumout;
wire fxp_functions_0_aadd_16_a12;
wire fxp_functions_0_aadd_21_a37_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_19_a32_cout;
wire fxp_functions_0_aadd_14_a6_sumout;
wire fxp_functions_0_aadd_14_a7;
wire fxp_functions_0_aadd_17_a27_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_15_a22_cout;
wire fxp_functions_0_aadd_12_a1_sumout;
wire fxp_functions_0_aadd_13_a17_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a8_a_aq;
wire fxp_functions_0_aadd_11_a12_cout;
wire fxp_functions_0_aadd_9_a7_cout;
wire fxp_functions_0_aadd_7_a1_sumout;
wire fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a_aq;
wire fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a_aq;
wire fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a_aq;
wire fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a_aq;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_20_a26_sumout;
wire fxp_functions_0_aadd_20_a27;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_22_a31_sumout;
wire fxp_functions_0_aadd_22_a32;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_24_a36_sumout;
wire fxp_functions_0_aadd_24_a37;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_26_a41_sumout;
wire fxp_functions_0_aadd_26_a42;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_28_a46_sumout;
wire fxp_functions_0_aadd_28_a47;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_29_a62_cout;
wire fxp_functions_0_aadd_30_a51_sumout;
wire fxp_functions_0_aadd_30_a52;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a7_a_aq;
wire fxp_functions_0_aadd_31_a67_cout;
wire fxp_functions_0_aadd_18_a21_sumout;
wire fxp_functions_0_aadd_18_a22;
wire fxp_functions_0_aadd_27_a57_cout;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_25_a52_cout;
wire fxp_functions_0_aadd_16_a16_sumout;
wire fxp_functions_0_aadd_16_a17;
wire fxp_functions_0_aadd_23_a47_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_21_a42_cout;
wire fxp_functions_0_aadd_14_a11_sumout;
wire fxp_functions_0_aadd_14_a12;
wire fxp_functions_0_aadd_19_a37_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_17_a32_cout;
wire fxp_functions_0_aadd_12_a6_sumout;
wire fxp_functions_0_aadd_12_a7;
wire fxp_functions_0_aadd_15_a27_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_13_a22_cout;
wire fxp_functions_0_aadd_10_a1_sumout;
wire fxp_functions_0_aadd_11_a17_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a7_a_aq;
wire fxp_functions_0_aadd_9_a12_cout;
wire fxp_functions_0_aadd_7_a7_cout;
wire fxp_functions_0_aadd_5_a1_sumout;
wire fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aadd_18_a26_sumout;
wire fxp_functions_0_aadd_18_a27;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_20_a31_sumout;
wire fxp_functions_0_aadd_20_a32;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_22_a36_sumout;
wire fxp_functions_0_aadd_22_a37;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_24_a41_sumout;
wire fxp_functions_0_aadd_24_a42;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_26_a46_sumout;
wire fxp_functions_0_aadd_26_a47;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_28_a51_sumout;
wire fxp_functions_0_aadd_28_a52;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_29_a67_cout;
wire fxp_functions_0_aadd_30_a56_sumout;
wire fxp_functions_0_aadd_30_a57;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a6_a_aq;
wire fxp_functions_0_aadd_31_a72_cout;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_27_a62_cout;
wire fxp_functions_0_aadd_16_a21_sumout;
wire fxp_functions_0_aadd_16_a22;
wire fxp_functions_0_aadd_25_a57_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_23_a52_cout;
wire fxp_functions_0_aadd_14_a16_sumout;
wire fxp_functions_0_aadd_14_a17;
wire fxp_functions_0_aadd_21_a47_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_19_a42_cout;
wire fxp_functions_0_aadd_12_a11_sumout;
wire fxp_functions_0_aadd_12_a12;
wire fxp_functions_0_aadd_17_a37_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_15_a32_cout;
wire fxp_functions_0_aadd_10_a6_sumout;
wire fxp_functions_0_aadd_10_a7;
wire fxp_functions_0_aadd_13_a27_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_11_a22_cout;
wire fxp_functions_0_aadd_8_a1_sumout;
wire fxp_functions_0_aadd_9_a17_cout;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a6_a_aq;
wire fxp_functions_0_aadd_7_a12_cout;
wire fxp_functions_0_aadd_5_a7_cout;
wire fxp_functions_0_aadd_3_a1_sumout;
wire fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq;
wire fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a_aq;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_18_a31_sumout;
wire fxp_functions_0_aadd_18_a32;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_20_a36_sumout;
wire fxp_functions_0_aadd_20_a37;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_22_a41_sumout;
wire fxp_functions_0_aadd_22_a42;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_24_a46_sumout;
wire fxp_functions_0_aadd_24_a47;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_26_a51_sumout;
wire fxp_functions_0_aadd_26_a52;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_28_a56_sumout;
wire fxp_functions_0_aadd_28_a57;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_29_a72_cout;
wire fxp_functions_0_aadd_30_a61_sumout;
wire fxp_functions_0_aadd_30_a62;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a5_a_aq;
wire fxp_functions_0_aadd_31_a77_cout;
wire fxp_functions_0_aadd_16_a26_sumout;
wire fxp_functions_0_aadd_16_a27;
wire fxp_functions_0_aadd_27_a67_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_25_a62_cout;
wire fxp_functions_0_aadd_14_a21_sumout;
wire fxp_functions_0_aadd_14_a22;
wire fxp_functions_0_aadd_23_a57_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_21_a52_cout;
wire fxp_functions_0_aadd_12_a16_sumout;
wire fxp_functions_0_aadd_12_a17;
wire fxp_functions_0_aadd_19_a47_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_17_a42_cout;
wire fxp_functions_0_aadd_10_a11_sumout;
wire fxp_functions_0_aadd_10_a12;
wire fxp_functions_0_aadd_15_a37_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_13_a32_cout;
wire fxp_functions_0_aadd_8_a6_sumout;
wire fxp_functions_0_aadd_8_a7;
wire fxp_functions_0_aadd_11_a27_cout;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_9_a22_cout;
wire fxp_functions_0_aadd_6_a1_sumout;
wire fxp_functions_0_aadd_7_a17_cout;
wire fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a5_a_aq;
wire fxp_functions_0_aadd_5_a12_cout;
wire fxp_functions_0_aadd_3_a7_cout;
wire fxp_functions_0_aadd_16_a31_sumout;
wire fxp_functions_0_aadd_16_a32;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_18_a36_sumout;
wire fxp_functions_0_aadd_18_a37;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_20_a41_sumout;
wire fxp_functions_0_aadd_20_a42;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_22_a46_sumout;
wire fxp_functions_0_aadd_22_a47;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_24_a51_sumout;
wire fxp_functions_0_aadd_24_a52;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_26_a56_sumout;
wire fxp_functions_0_aadd_26_a57;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_28_a61_sumout;
wire fxp_functions_0_aadd_28_a62;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_29_a77_cout;
wire fxp_functions_0_aadd_30_a66_sumout;
wire fxp_functions_0_aadd_30_a67;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a4_a_aq;
wire fxp_functions_0_aadd_31_a82_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_27_a72_cout;
wire fxp_functions_0_aadd_14_a26_sumout;
wire fxp_functions_0_aadd_14_a27;
wire fxp_functions_0_aadd_25_a67_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_23_a62_cout;
wire fxp_functions_0_aadd_12_a21_sumout;
wire fxp_functions_0_aadd_12_a22;
wire fxp_functions_0_aadd_21_a57_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_19_a52_cout;
wire fxp_functions_0_aadd_10_a16_sumout;
wire fxp_functions_0_aadd_10_a17;
wire fxp_functions_0_aadd_17_a47_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_15_a42_cout;
wire fxp_functions_0_aadd_8_a11_sumout;
wire fxp_functions_0_aadd_8_a12;
wire fxp_functions_0_aadd_13_a37_cout;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_11_a32_cout;
wire fxp_functions_0_aadd_6_a6_sumout;
wire fxp_functions_0_aadd_6_a7;
wire fxp_functions_0_aadd_9_a27_cout;
wire fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a_aq;
wire fxp_functions_0_aadd_7_a22_cout;
wire fxp_functions_0_aadd_4_a1_sumout;
wire fxp_functions_0_aadd_5_a17_cout;
wire fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_3_a12_cout;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_16_a36_sumout;
wire fxp_functions_0_aadd_16_a37;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_18_a41_sumout;
wire fxp_functions_0_aadd_18_a42;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_20_a46_sumout;
wire fxp_functions_0_aadd_20_a47;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_22_a51_sumout;
wire fxp_functions_0_aadd_22_a52;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_24_a56_sumout;
wire fxp_functions_0_aadd_24_a57;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_26_a61_sumout;
wire fxp_functions_0_aadd_26_a62;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_28_a66_sumout;
wire fxp_functions_0_aadd_28_a67;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_29_a82_cout;
wire fxp_functions_0_aadd_30_a71_sumout;
wire fxp_functions_0_aadd_30_a72;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a3_a_aq;
wire fxp_functions_0_aadd_31_a87_cout;
wire fxp_functions_0_aadd_14_a31_sumout;
wire fxp_functions_0_aadd_14_a32;
wire fxp_functions_0_aadd_27_a77_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_25_a72_cout;
wire fxp_functions_0_aadd_12_a26_sumout;
wire fxp_functions_0_aadd_12_a27;
wire fxp_functions_0_aadd_23_a67_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_21_a62_cout;
wire fxp_functions_0_aadd_10_a21_sumout;
wire fxp_functions_0_aadd_10_a22;
wire fxp_functions_0_aadd_19_a57_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_17_a52_cout;
wire fxp_functions_0_aadd_8_a16_sumout;
wire fxp_functions_0_aadd_8_a17;
wire fxp_functions_0_aadd_15_a47_cout;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_13_a42_cout;
wire fxp_functions_0_aadd_6_a11_sumout;
wire fxp_functions_0_aadd_6_a12;
wire fxp_functions_0_aadd_11_a37_cout;
wire fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a_aq;
wire fxp_functions_0_aadd_9_a32_cout;
wire fxp_functions_0_aadd_4_a6_sumout;
wire fxp_functions_0_aadd_4_a7;
wire fxp_functions_0_aadd_7_a27_cout;
wire fxp_functions_0_aadd_5_a22_cout;
wire fxp_functions_0_aadd_3_a17_cout;
wire fxp_functions_0_aadd_14_a36_sumout;
wire fxp_functions_0_aadd_14_a37;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_16_a41_sumout;
wire fxp_functions_0_aadd_16_a42;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_18_a46_sumout;
wire fxp_functions_0_aadd_18_a47;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_20_a51_sumout;
wire fxp_functions_0_aadd_20_a52;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_22_a56_sumout;
wire fxp_functions_0_aadd_22_a57;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_24_a61_sumout;
wire fxp_functions_0_aadd_24_a62;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_26_a66_sumout;
wire fxp_functions_0_aadd_26_a67;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_28_a71_sumout;
wire fxp_functions_0_aadd_28_a72;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_29_a87_cout;
wire fxp_functions_0_aadd_30_a76_sumout;
wire fxp_functions_0_aadd_30_a77;
wire fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_27_a82_cout;
wire fxp_functions_0_aadd_12_a31_sumout;
wire fxp_functions_0_aadd_12_a32;
wire fxp_functions_0_aadd_25_a77_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_23_a72_cout;
wire fxp_functions_0_aadd_10_a26_sumout;
wire fxp_functions_0_aadd_10_a27;
wire fxp_functions_0_aadd_21_a67_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_19_a62_cout;
wire fxp_functions_0_aadd_8_a21_sumout;
wire fxp_functions_0_aadd_8_a22;
wire fxp_functions_0_aadd_17_a57_cout;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_15_a52_cout;
wire fxp_functions_0_aadd_6_a16_sumout;
wire fxp_functions_0_aadd_6_a17;
wire fxp_functions_0_aadd_13_a47_cout;
wire fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a_aq;
wire fxp_functions_0_aadd_11_a42_cout;
wire fxp_functions_0_aadd_4_a11_sumout;
wire fxp_functions_0_aadd_4_a12;
wire fxp_functions_0_aadd_9_a37_cout;
wire fxp_functions_0_aadd_7_a32_cout;
wire fxp_functions_0_aadd_5_a27_cout;
wire fxp_functions_0_aadd_3_a22_cout;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_14_a41_sumout;
wire fxp_functions_0_aadd_14_a42;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_16_a46_sumout;
wire fxp_functions_0_aadd_16_a47;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_18_a51_sumout;
wire fxp_functions_0_aadd_18_a52;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_20_a56_sumout;
wire fxp_functions_0_aadd_20_a57;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_22_a61_sumout;
wire fxp_functions_0_aadd_22_a62;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_24_a66_sumout;
wire fxp_functions_0_aadd_24_a67;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_26_a71_sumout;
wire fxp_functions_0_aadd_26_a72;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_28_a76_sumout;
wire fxp_functions_0_aadd_28_a77;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_29_a92_cout;
wire fxp_functions_0_aadd_30_a81_sumout;
wire fxp_functions_0_aadd_30_a82;
wire fxp_functions_0_aadd_12_a36_sumout;
wire fxp_functions_0_aadd_12_a37;
wire fxp_functions_0_aadd_27_a87_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_25_a82_cout;
wire fxp_functions_0_aadd_10_a31_sumout;
wire fxp_functions_0_aadd_10_a32;
wire fxp_functions_0_aadd_23_a77_cout;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_21_a72_cout;
wire fxp_functions_0_aadd_8_a26_sumout;
wire fxp_functions_0_aadd_8_a27;
wire fxp_functions_0_aadd_19_a67_cout;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_17_a62_cout;
wire fxp_functions_0_aadd_6_a21_sumout;
wire fxp_functions_0_aadd_6_a22;
wire fxp_functions_0_aadd_15_a57_cout;
wire fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a_aq;
wire fxp_functions_0_aadd_13_a52_cout;
wire fxp_functions_0_aadd_4_a16_sumout;
wire fxp_functions_0_aadd_4_a17;
wire fxp_functions_0_aadd_11_a47_cout;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a_aq;
wire fxp_functions_0_aadd_9_a42_cout;
wire fxp_functions_0_aadd_7_a37_cout;
wire fxp_functions_0_aadd_5_a32_cout;
wire fxp_functions_0_aadd_3_a27_cout;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_14_a47_cout;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_16_a52_cout;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_18_a57_cout;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_20_a62_cout;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_22_a67_cout;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_24_a72_cout;
wire fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_26_a77_cout;
wire fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_28_a82_cout;
wire fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_30_a87_cout;
wire fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_12_a42_cout;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_10_a37_cout;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a23_a_aq;
wire fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_8_a32_cout;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a25_a_aq;
wire fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a_aq;
wire fxp_functions_0_aadd_6_a27_cout;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a27_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a_aq;
wire fxp_functions_0_aadd_4_a22_cout;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a22_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a23_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a24_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a25_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a26_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a22_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a23_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a24_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a22_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout;
wire fxp_functions_0_aadd_1_a0_combout;
wire fxp_functions_0_areduce_nor_0_acombout;
wire fxp_functions_0_aadd_2_a0_combout;
wire fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0_combout;
wire fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0_combout;
wire fxp_functions_0_ai240_a0_combout;
wire fxp_functions_0_aadd_0_a0_combout;
wire a_aGND_acombout;
wire fxp_functions_0_aadd_11_a1_wirecell_combout;
wire fxp_functions_0_aadd_13_a1_wirecell_combout;
wire fxp_functions_0_aadd_15_a1_wirecell_combout;
wire fxp_functions_0_aadd_17_a1_wirecell_combout;
wire fxp_functions_0_aadd_19_a1_wirecell_combout;
wire fxp_functions_0_aadd_21_a1_wirecell_combout;
wire fxp_functions_0_aadd_23_a1_wirecell_combout;
wire fxp_functions_0_aadd_25_a1_wirecell_combout;
wire fxp_functions_0_aadd_27_a1_wirecell_combout;
wire fxp_functions_0_aadd_29_a1_wirecell_combout;
wire fxp_functions_0_aadd_3_a1_wirecell_combout;
wire fxp_functions_0_aadd_5_a1_wirecell_combout;
wire fxp_functions_0_aadd_7_a1_wirecell_combout;
wire fxp_functions_0_aadd_9_a1_wirecell_combout;
wire fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell_combout;


fourteennm_lcell_comb fxp_functions_0_aadd_32_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_31_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a1_sumout),
	.cout(fxp_functions_0_aadd_32_a2),
	.shareout());
defparam fxp_functions_0_aadd_32_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a1.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_32_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a6_sumout),
	.cout(fxp_functions_0_aadd_32_a7),
	.shareout());
defparam fxp_functions_0_aadd_32_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a6.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a11_sumout),
	.cout(fxp_functions_0_aadd_32_a12),
	.shareout());
defparam fxp_functions_0_aadd_32_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a11.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a16_sumout),
	.cout(fxp_functions_0_aadd_32_a17),
	.shareout());
defparam fxp_functions_0_aadd_32_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a16.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a21_sumout),
	.cout(fxp_functions_0_aadd_32_a22),
	.shareout());
defparam fxp_functions_0_aadd_32_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a21.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a26_sumout),
	.cout(fxp_functions_0_aadd_32_a27),
	.shareout());
defparam fxp_functions_0_aadd_32_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a26.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a31_sumout),
	.cout(fxp_functions_0_aadd_32_a32),
	.shareout());
defparam fxp_functions_0_aadd_32_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a31.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a36_sumout),
	.cout(fxp_functions_0_aadd_32_a37),
	.shareout());
defparam fxp_functions_0_aadd_32_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a36.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a41_sumout),
	.cout(fxp_functions_0_aadd_32_a42),
	.shareout());
defparam fxp_functions_0_aadd_32_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a41.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a46_sumout),
	.cout(fxp_functions_0_aadd_32_a47),
	.shareout());
defparam fxp_functions_0_aadd_32_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a46.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a51_sumout),
	.cout(fxp_functions_0_aadd_32_a52),
	.shareout());
defparam fxp_functions_0_aadd_32_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a51.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a56_sumout),
	.cout(fxp_functions_0_aadd_32_a57),
	.shareout());
defparam fxp_functions_0_aadd_32_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a56.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a61_sumout),
	.cout(fxp_functions_0_aadd_32_a62),
	.shareout());
defparam fxp_functions_0_aadd_32_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a61.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a66_sumout),
	.cout(fxp_functions_0_aadd_32_a67),
	.shareout());
defparam fxp_functions_0_aadd_32_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a66.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a71_sumout),
	.cout(fxp_functions_0_aadd_32_a72),
	.shareout());
defparam fxp_functions_0_aadd_32_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a71.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a76_sumout),
	.cout(fxp_functions_0_aadd_32_a77),
	.shareout());
defparam fxp_functions_0_aadd_32_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a76.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_32_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_32_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_32_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_32_a81_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_32_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_32_a81.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_aadd_32_a81.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_29_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_31_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_31_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_31_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a_aq));
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_29_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_29_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_29_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_31_a7.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_27_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a_aq));
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_29_a7.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a18_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a15_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a17_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_27_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_27_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_27_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_25_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a_aq));
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a17_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a1(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a14_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_30_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_30_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a14_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a16_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_27_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_25_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_25_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_25_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_23_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a_aq));
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a1(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_28_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_28_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a16_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a17.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a6(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a13_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a6_sumout),
	.cout(fxp_functions_0_aadd_30_a7),
	.shareout());
defparam fxp_functions_0_aadd_30_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a6.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a16_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a15_a_aq),
	.datad(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a22.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_31_a22.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a16_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a16_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_25_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_23_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_23_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_23_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_21_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a_aq));
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a6(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a6_sumout),
	.cout(fxp_functions_0_aadd_28_a7),
	.shareout());
defparam fxp_functions_0_aadd_28_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a6.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a22.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a11(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a11_sumout),
	.cout(fxp_functions_0_aadd_30_a12),
	.shareout());
defparam fxp_functions_0_aadd_30_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a11.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a14_a_aq),
	.datad(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a27.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_31_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a1(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_26_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_26_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a17.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a15_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_23_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_21_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_21_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_21_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_19_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a_aq));
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a6(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a6_sumout),
	.cout(fxp_functions_0_aadd_26_a7),
	.shareout());
defparam fxp_functions_0_aadd_26_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a6.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a14_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a11(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a11_sumout),
	.cout(fxp_functions_0_aadd_28_a12),
	.shareout());
defparam fxp_functions_0_aadd_28_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a11.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a14_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a27.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a16(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a16_sumout),
	.cout(fxp_functions_0_aadd_30_a17),
	.shareout());
defparam fxp_functions_0_aadd_30_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a16.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a14_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a13_a_aq),
	.datad(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a32.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_31_a32.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a14_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a22.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a1(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_24_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_24_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a14_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a14_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_21_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_19_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_19_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_19_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a_aq));
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a11(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a11_sumout),
	.cout(fxp_functions_0_aadd_26_a12),
	.shareout());
defparam fxp_functions_0_aadd_26_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a11.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a16(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a16_sumout),
	.cout(fxp_functions_0_aadd_28_a17),
	.shareout());
defparam fxp_functions_0_aadd_28_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a16.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a32.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a21(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a21_sumout),
	.cout(fxp_functions_0_aadd_30_a22),
	.shareout());
defparam fxp_functions_0_aadd_30_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a37.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a6(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a6_sumout),
	.cout(fxp_functions_0_aadd_24_a7),
	.shareout());
defparam fxp_functions_0_aadd_24_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a27.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a1(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_22_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_22_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a13_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_21_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_19_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_17_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_17_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_15_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a_aq));
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a11(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a11_sumout),
	.cout(fxp_functions_0_aadd_24_a12),
	.shareout());
defparam fxp_functions_0_aadd_24_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a11.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a16(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a16_sumout),
	.cout(fxp_functions_0_aadd_26_a17),
	.shareout());
defparam fxp_functions_0_aadd_26_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a16.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a21(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a21_sumout),
	.cout(fxp_functions_0_aadd_28_a22),
	.shareout());
defparam fxp_functions_0_aadd_28_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a37.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a37.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a26(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a26_sumout),
	.cout(fxp_functions_0_aadd_30_a27),
	.shareout());
defparam fxp_functions_0_aadd_30_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a42.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_31_a42.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a32.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a6(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a6_sumout),
	.cout(fxp_functions_0_aadd_22_a7),
	.shareout());
defparam fxp_functions_0_aadd_22_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a1(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_20_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_20_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a17.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_21_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a12_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a12_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datad(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_19_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_17_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_15_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_15_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_15_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a_aq));
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a16(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a16_sumout),
	.cout(fxp_functions_0_aadd_24_a17),
	.shareout());
defparam fxp_functions_0_aadd_24_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a16.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a21(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a21_sumout),
	.cout(fxp_functions_0_aadd_26_a22),
	.shareout());
defparam fxp_functions_0_aadd_26_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a26(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a26_sumout),
	.cout(fxp_functions_0_aadd_28_a27),
	.shareout());
defparam fxp_functions_0_aadd_28_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a42.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a31(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a31_sumout),
	.cout(fxp_functions_0_aadd_30_a32),
	.shareout());
defparam fxp_functions_0_aadd_30_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a47.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a47.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a11(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a11_sumout),
	.cout(fxp_functions_0_aadd_22_a12),
	.shareout());
defparam fxp_functions_0_aadd_22_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a37.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a6(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a6_sumout),
	.cout(fxp_functions_0_aadd_20_a7),
	.shareout());
defparam fxp_functions_0_aadd_20_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a22.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_21_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a1(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_18_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_18_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a17.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_19_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a11_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_17_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_15_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_13_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_13_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_11_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a_aq));
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a16(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a16_sumout),
	.cout(fxp_functions_0_aadd_22_a17),
	.shareout());
defparam fxp_functions_0_aadd_22_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a16.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a21(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a21_sumout),
	.cout(fxp_functions_0_aadd_24_a22),
	.shareout());
defparam fxp_functions_0_aadd_24_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a26(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a26_sumout),
	.cout(fxp_functions_0_aadd_26_a27),
	.shareout());
defparam fxp_functions_0_aadd_26_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a31(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a31_sumout),
	.cout(fxp_functions_0_aadd_28_a32),
	.shareout());
defparam fxp_functions_0_aadd_28_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a47.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a47.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a36(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a36_sumout),
	.cout(fxp_functions_0_aadd_30_a37),
	.shareout());
defparam fxp_functions_0_aadd_30_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a52.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a52.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a42.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a11(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a11_sumout),
	.cout(fxp_functions_0_aadd_20_a12),
	.shareout());
defparam fxp_functions_0_aadd_20_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a6(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a6_sumout),
	.cout(fxp_functions_0_aadd_18_a7),
	.shareout());
defparam fxp_functions_0_aadd_18_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a22.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_19_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a1(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_16_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_16_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a10_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_15_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_13_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_11_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_11_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_11_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a21(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a21_sumout),
	.cout(fxp_functions_0_aadd_22_a22),
	.shareout());
defparam fxp_functions_0_aadd_22_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a26(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a26_sumout),
	.cout(fxp_functions_0_aadd_24_a27),
	.shareout());
defparam fxp_functions_0_aadd_24_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a31(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a31_sumout),
	.cout(fxp_functions_0_aadd_26_a32),
	.shareout());
defparam fxp_functions_0_aadd_26_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a36(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a36_sumout),
	.cout(fxp_functions_0_aadd_28_a37),
	.shareout());
defparam fxp_functions_0_aadd_28_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a52.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a41(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a41_sumout),
	.cout(fxp_functions_0_aadd_30_a42),
	.shareout());
defparam fxp_functions_0_aadd_30_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a57.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a57.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a16(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a16_sumout),
	.cout(fxp_functions_0_aadd_20_a17),
	.shareout());
defparam fxp_functions_0_aadd_20_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a47.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a42.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a11(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a11_sumout),
	.cout(fxp_functions_0_aadd_18_a12),
	.shareout());
defparam fxp_functions_0_aadd_18_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a6(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a6_sumout),
	.cout(fxp_functions_0_aadd_16_a7),
	.shareout());
defparam fxp_functions_0_aadd_16_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a1(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_14_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_14_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_15_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a9_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_13_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_11_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_9_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_9_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a21(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a21_sumout),
	.cout(fxp_functions_0_aadd_20_a22),
	.shareout());
defparam fxp_functions_0_aadd_20_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a26(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a26_sumout),
	.cout(fxp_functions_0_aadd_22_a27),
	.shareout());
defparam fxp_functions_0_aadd_22_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a31(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a31_sumout),
	.cout(fxp_functions_0_aadd_24_a32),
	.shareout());
defparam fxp_functions_0_aadd_24_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a36(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a36_sumout),
	.cout(fxp_functions_0_aadd_26_a37),
	.shareout());
defparam fxp_functions_0_aadd_26_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a41(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a41_sumout),
	.cout(fxp_functions_0_aadd_28_a42),
	.shareout());
defparam fxp_functions_0_aadd_28_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a57.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a57.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a46(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a46_sumout),
	.cout(fxp_functions_0_aadd_30_a47),
	.shareout());
defparam fxp_functions_0_aadd_30_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a46.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a62.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a62.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a52.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a16(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a16_sumout),
	.cout(fxp_functions_0_aadd_18_a17),
	.shareout());
defparam fxp_functions_0_aadd_18_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a47.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a42.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_23_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a11(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a11_sumout),
	.cout(fxp_functions_0_aadd_16_a12),
	.shareout());
defparam fxp_functions_0_aadd_16_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a6(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a6_sumout),
	.cout(fxp_functions_0_aadd_14_a7),
	.shareout());
defparam fxp_functions_0_aadd_14_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_14_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_15_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a1(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_12_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_12_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_13_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a8_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_11_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_9_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_7_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_7_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_5_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a_aq));
defparam fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a_aq));
defparam fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a_aq));
defparam fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a_aq));
defparam fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a26(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a26_sumout),
	.cout(fxp_functions_0_aadd_20_a27),
	.shareout());
defparam fxp_functions_0_aadd_20_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a31(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a31_sumout),
	.cout(fxp_functions_0_aadd_22_a32),
	.shareout());
defparam fxp_functions_0_aadd_22_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a36(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a36_sumout),
	.cout(fxp_functions_0_aadd_24_a37),
	.shareout());
defparam fxp_functions_0_aadd_24_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a41(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a41_sumout),
	.cout(fxp_functions_0_aadd_26_a42),
	.shareout());
defparam fxp_functions_0_aadd_26_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a46(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a46_sumout),
	.cout(fxp_functions_0_aadd_28_a47),
	.shareout());
defparam fxp_functions_0_aadd_28_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a46.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a62.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_29_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a51(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a51_sumout),
	.cout(fxp_functions_0_aadd_30_a52),
	.shareout());
defparam fxp_functions_0_aadd_30_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a51.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a67.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a67.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a21(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a21_sumout),
	.cout(fxp_functions_0_aadd_18_a22),
	.shareout());
defparam fxp_functions_0_aadd_18_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a57.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a52.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a16(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a16_sumout),
	.cout(fxp_functions_0_aadd_16_a17),
	.shareout());
defparam fxp_functions_0_aadd_16_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a47.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_23_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a42.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a11(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a11_sumout),
	.cout(fxp_functions_0_aadd_14_a12),
	.shareout());
defparam fxp_functions_0_aadd_14_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_14_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a6(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a6_sumout),
	.cout(fxp_functions_0_aadd_12_a7),
	.shareout());
defparam fxp_functions_0_aadd_12_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_12_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_15_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_13_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a1(
	.dataa(!fxp_functions_0_aadd_9_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_10_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_10_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_11_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a7_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_9_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_7_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_5_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_5_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_5_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_5_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_3_a1_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a26(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a26_sumout),
	.cout(fxp_functions_0_aadd_18_a27),
	.shareout());
defparam fxp_functions_0_aadd_18_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a26.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a31(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a31_sumout),
	.cout(fxp_functions_0_aadd_20_a32),
	.shareout());
defparam fxp_functions_0_aadd_20_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a36(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a36_sumout),
	.cout(fxp_functions_0_aadd_22_a37),
	.shareout());
defparam fxp_functions_0_aadd_22_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a41(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a41_sumout),
	.cout(fxp_functions_0_aadd_24_a42),
	.shareout());
defparam fxp_functions_0_aadd_24_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a46(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a46_sumout),
	.cout(fxp_functions_0_aadd_26_a47),
	.shareout());
defparam fxp_functions_0_aadd_26_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a46.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a51(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a51_sumout),
	.cout(fxp_functions_0_aadd_28_a52),
	.shareout());
defparam fxp_functions_0_aadd_28_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a51.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a67.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_29_a67.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a56(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a56_sumout),
	.cout(fxp_functions_0_aadd_30_a57),
	.shareout());
defparam fxp_functions_0_aadd_30_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a56.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a56.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a72.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a72.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a62.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a21(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a21_sumout),
	.cout(fxp_functions_0_aadd_16_a22),
	.shareout());
defparam fxp_functions_0_aadd_16_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a57.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a52.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_23_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a16(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a16_sumout),
	.cout(fxp_functions_0_aadd_14_a17),
	.shareout());
defparam fxp_functions_0_aadd_14_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_14_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a47.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a42.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a11(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a11_sumout),
	.cout(fxp_functions_0_aadd_12_a12),
	.shareout());
defparam fxp_functions_0_aadd_12_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_12_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_15_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a6(
	.dataa(!fxp_functions_0_aadd_9_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a6_sumout),
	.cout(fxp_functions_0_aadd_10_a7),
	.shareout());
defparam fxp_functions_0_aadd_10_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_10_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_13_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_11_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a1(
	.dataa(!fxp_functions_0_aadd_7_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_8_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_8_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_9_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_6_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a6_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a12.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_7_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_5_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_5_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_5_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_5_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_3_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_3_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_3_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a1.lut_mask = 64'h000000000000FFFF;
defparam fxp_functions_0_aadd_3_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_1_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq));
defparam fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_0_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a31(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a31_sumout),
	.cout(fxp_functions_0_aadd_18_a32),
	.shareout());
defparam fxp_functions_0_aadd_18_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a36(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a36_sumout),
	.cout(fxp_functions_0_aadd_20_a37),
	.shareout());
defparam fxp_functions_0_aadd_20_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a41(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a41_sumout),
	.cout(fxp_functions_0_aadd_22_a42),
	.shareout());
defparam fxp_functions_0_aadd_22_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a46(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a46_sumout),
	.cout(fxp_functions_0_aadd_24_a47),
	.shareout());
defparam fxp_functions_0_aadd_24_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a46.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a51(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a51_sumout),
	.cout(fxp_functions_0_aadd_26_a52),
	.shareout());
defparam fxp_functions_0_aadd_26_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a51.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a56(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a56_sumout),
	.cout(fxp_functions_0_aadd_28_a57),
	.shareout());
defparam fxp_functions_0_aadd_28_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a56.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a56.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a72.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_29_a72.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a61(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a61_sumout),
	.cout(fxp_functions_0_aadd_30_a62),
	.shareout());
defparam fxp_functions_0_aadd_30_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a61.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a61.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a82_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a77_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a77.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a77.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a77.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a26(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a26_sumout),
	.cout(fxp_functions_0_aadd_16_a27),
	.shareout());
defparam fxp_functions_0_aadd_16_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a67.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a67.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a62.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a21(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a21_sumout),
	.cout(fxp_functions_0_aadd_14_a22),
	.shareout());
defparam fxp_functions_0_aadd_14_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_14_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a57.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a52.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a16(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a16_sumout),
	.cout(fxp_functions_0_aadd_12_a17),
	.shareout());
defparam fxp_functions_0_aadd_12_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_12_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a47.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a42.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a11(
	.dataa(!fxp_functions_0_aadd_9_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a11_sumout),
	.cout(fxp_functions_0_aadd_10_a12),
	.shareout());
defparam fxp_functions_0_aadd_10_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_10_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_15_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a32.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_13_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a6(
	.dataa(!fxp_functions_0_aadd_7_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a6_sumout),
	.cout(fxp_functions_0_aadd_8_a7),
	.shareout());
defparam fxp_functions_0_aadd_8_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_8_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_11_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_6_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_9_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_6_a1(
	.dataa(!fxp_functions_0_aadd_5_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_6_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_6_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_6_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_6_a1.lut_mask = 64'h000000000000F50A;
defparam fxp_functions_0_aadd_6_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a17.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_7_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_4_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a5_a_aq));
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_5_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_5_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_5_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a12.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_5_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aadd_2_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_3_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_3_a7_cout),
	.shareout());
defparam fxp_functions_0_aadd_3_a7.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a7.lut_mask = 64'h00000000F0F00F0F;
defparam fxp_functions_0_aadd_3_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a31(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a31_sumout),
	.cout(fxp_functions_0_aadd_16_a32),
	.shareout());
defparam fxp_functions_0_aadd_16_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a31.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a36(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a36_sumout),
	.cout(fxp_functions_0_aadd_18_a37),
	.shareout());
defparam fxp_functions_0_aadd_18_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a41(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a41_sumout),
	.cout(fxp_functions_0_aadd_20_a42),
	.shareout());
defparam fxp_functions_0_aadd_20_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a46(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a46_sumout),
	.cout(fxp_functions_0_aadd_22_a47),
	.shareout());
defparam fxp_functions_0_aadd_22_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a46.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a51(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a51_sumout),
	.cout(fxp_functions_0_aadd_24_a52),
	.shareout());
defparam fxp_functions_0_aadd_24_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a51.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a56(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a56_sumout),
	.cout(fxp_functions_0_aadd_26_a57),
	.shareout());
defparam fxp_functions_0_aadd_26_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a56.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a56.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a61(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a61_sumout),
	.cout(fxp_functions_0_aadd_28_a62),
	.shareout());
defparam fxp_functions_0_aadd_28_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a61.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a61.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a82_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a77_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a77.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a77.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_29_a77.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a66(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a66_sumout),
	.cout(fxp_functions_0_aadd_30_a67),
	.shareout());
defparam fxp_functions_0_aadd_30_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a66.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a66.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a82(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_31_a87_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a82_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a82.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a82.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a82.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a72.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a72.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a26(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a26_sumout),
	.cout(fxp_functions_0_aadd_14_a27),
	.shareout());
defparam fxp_functions_0_aadd_14_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_14_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a67.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a67.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a62.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_23_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a21(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a21_sumout),
	.cout(fxp_functions_0_aadd_12_a22),
	.shareout());
defparam fxp_functions_0_aadd_12_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_12_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a57.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a52.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a16(
	.dataa(!fxp_functions_0_aadd_9_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a16_sumout),
	.cout(fxp_functions_0_aadd_10_a17),
	.shareout());
defparam fxp_functions_0_aadd_10_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_10_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a47.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a42.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_15_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a11(
	.dataa(!fxp_functions_0_aadd_7_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a11_sumout),
	.cout(fxp_functions_0_aadd_8_a12),
	.shareout());
defparam fxp_functions_0_aadd_8_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_8_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_13_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_6_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_11_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_6_a6(
	.dataa(!fxp_functions_0_aadd_5_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_6_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_6_a6_sumout),
	.cout(fxp_functions_0_aadd_6_a7),
	.shareout());
defparam fxp_functions_0_aadd_6_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_6_a6.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_6_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a27.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_9_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_4_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a_aq));
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist43_sM_plus2pow_uid38_sqrt_q_2_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a22.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_7_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_4_a1(
	.dataa(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datab(!fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0_combout),
	.datac(!fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0_combout),
	.datad(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_4_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_4_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_4_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_4_a1.lut_mask = 64'h000000000000D22D;
defparam fxp_functions_0_aadd_4_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_5_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_5_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_5_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a17.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_5_a17.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai240_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(radical[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(radical[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_0_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a12(
	.dataa(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datab(!fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0_combout),
	.datac(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_3_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_3_a12_cout),
	.shareout());
defparam fxp_functions_0_aadd_3_a12.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a12.lut_mask = 64'h000000002D00D22D;
defparam fxp_functions_0_aadd_3_a12.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a36(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a36_sumout),
	.cout(fxp_functions_0_aadd_16_a37),
	.shareout());
defparam fxp_functions_0_aadd_16_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a36.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_16_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a41(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a41_sumout),
	.cout(fxp_functions_0_aadd_18_a42),
	.shareout());
defparam fxp_functions_0_aadd_18_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a41.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_18_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a46(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a46_sumout),
	.cout(fxp_functions_0_aadd_20_a47),
	.shareout());
defparam fxp_functions_0_aadd_20_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a46.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_20_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a51(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a51_sumout),
	.cout(fxp_functions_0_aadd_22_a52),
	.shareout());
defparam fxp_functions_0_aadd_22_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a51.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_22_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a56(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a56_sumout),
	.cout(fxp_functions_0_aadd_24_a57),
	.shareout());
defparam fxp_functions_0_aadd_24_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a56.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_24_a56.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a61(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a61_sumout),
	.cout(fxp_functions_0_aadd_26_a62),
	.shareout());
defparam fxp_functions_0_aadd_26_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a61.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_26_a61.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a66(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a66_sumout),
	.cout(fxp_functions_0_aadd_28_a67),
	.shareout());
defparam fxp_functions_0_aadd_28_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a66.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_28_a66.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a82(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a87_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a82_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a82.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a82.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_29_a82.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a71(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist30_sM_plus2pow_uid158_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a71_sumout),
	.cout(fxp_functions_0_aadd_30_a72),
	.shareout());
defparam fxp_functions_0_aadd_30_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a71.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_30_a71.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_31_a87(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist29_sM_plus2pow_uid168_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_31_a87_cout),
	.shareout());
defparam fxp_functions_0_aadd_31_a87.extended_lut = "off";
defparam fxp_functions_0_aadd_31_a87.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_31_a87.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a31(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a31_sumout),
	.cout(fxp_functions_0_aadd_14_a32),
	.shareout());
defparam fxp_functions_0_aadd_14_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a31.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_14_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist31_sM_plus2pow_uid148_sqrt_q_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a82_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a77_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a77.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a77.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_27_a77.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist32_sM_plus2pow_uid138_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a72.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_25_a72.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a26(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a26_sumout),
	.cout(fxp_functions_0_aadd_12_a27),
	.shareout());
defparam fxp_functions_0_aadd_12_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a26.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_12_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist33_sM_plus2pow_uid128_sqrt_q_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a67.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_23_a67.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist34_sM_plus2pow_uid118_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a62.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_21_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a21(
	.dataa(!fxp_functions_0_aadd_9_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a21_sumout),
	.cout(fxp_functions_0_aadd_10_a22),
	.shareout());
defparam fxp_functions_0_aadd_10_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a21.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_10_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist35_sM_plus2pow_uid108_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a57.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_19_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist36_sM_plus2pow_uid98_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a52.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_17_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a16(
	.dataa(!fxp_functions_0_aadd_7_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a16_sumout),
	.cout(fxp_functions_0_aadd_8_a17),
	.shareout());
defparam fxp_functions_0_aadd_8_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a16.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_8_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist37_sM_plus2pow_uid88_sqrt_q_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a47.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_15_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_6_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist38_sM_plus2pow_uid78_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a42.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_13_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_6_a11(
	.dataa(!fxp_functions_0_aadd_5_a1_sumout),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_6_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_6_a11_sumout),
	.cout(fxp_functions_0_aadd_6_a12),
	.shareout());
defparam fxp_functions_0_aadd_6_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_6_a11.lut_mask = 64'h0000000000F5F50A;
defparam fxp_functions_0_aadd_6_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist39_sM_plus2pow_uid68_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a37.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_11_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_4_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a_aq));
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist40_sM_plus2pow_uid58_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a32.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_9_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_4_a6(
	.dataa(!fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq),
	.datab(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aadd_3_a1_sumout),
	.datad(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_4_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_4_a6_sumout),
	.cout(fxp_functions_0_aadd_4_a7),
	.shareout());
defparam fxp_functions_0_aadd_4_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_4_a6.lut_mask = 64'h0000000013196CC6;
defparam fxp_functions_0_aadd_4_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist41_sE_cmpge_uid43_sqrt_n_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a27.lut_mask = 64'h000000000F00F00F;
defparam fxp_functions_0_aadd_7_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist42_sM_plus2pow_uid38_sqrt_q_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_5_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_5_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_5_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a22.lut_mask = 64'h0000000000F0F00F;
defparam fxp_functions_0_aadd_5_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a17(
	.dataa(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datab(!fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0_combout),
	.datac(gnd),
	.datad(!fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_3_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_3_a17_cout),
	.shareout());
defparam fxp_functions_0_aadd_3_a17.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a17.lut_mask = 64'h0000000000666699;
defparam fxp_functions_0_aadd_3_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a36_sumout),
	.cout(fxp_functions_0_aadd_14_a37),
	.shareout());
defparam fxp_functions_0_aadd_14_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a36.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_14_a36.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_14_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a41_sumout),
	.cout(fxp_functions_0_aadd_16_a42),
	.shareout());
defparam fxp_functions_0_aadd_16_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a41.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_16_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_16_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a46_sumout),
	.cout(fxp_functions_0_aadd_18_a47),
	.shareout());
defparam fxp_functions_0_aadd_18_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a46.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_18_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_18_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a51_sumout),
	.cout(fxp_functions_0_aadd_20_a52),
	.shareout());
defparam fxp_functions_0_aadd_20_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a51.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_20_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_20_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a56_sumout),
	.cout(fxp_functions_0_aadd_22_a57),
	.shareout());
defparam fxp_functions_0_aadd_22_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a56.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_22_a56.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_22_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a61_sumout),
	.cout(fxp_functions_0_aadd_24_a62),
	.shareout());
defparam fxp_functions_0_aadd_24_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a61.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_24_a61.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_24_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a66_sumout),
	.cout(fxp_functions_0_aadd_26_a67),
	.shareout());
defparam fxp_functions_0_aadd_26_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a66.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_26_a66.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_26_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a71_sumout),
	.cout(fxp_functions_0_aadd_28_a72),
	.shareout());
defparam fxp_functions_0_aadd_28_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a71.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_28_a71.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_28_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a87(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_29_a92_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a87_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a87.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a87.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_29_a87.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a76_sumout),
	.cout(fxp_functions_0_aadd_30_a77),
	.shareout());
defparam fxp_functions_0_aadd_30_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a76.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_30_a76.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_30_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist28_sE_opinls_uid171_sqrt_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_12_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a82(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_27_a87_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a82_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a82.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a82.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_27_a82.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a31_sumout),
	.cout(fxp_functions_0_aadd_12_a32),
	.shareout());
defparam fxp_functions_0_aadd_12_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a31.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_12_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_25_a82_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a77_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a77.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a77.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_25_a77.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_10_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_23_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a72.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_23_a72.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a26_sumout),
	.cout(fxp_functions_0_aadd_10_a27),
	.shareout());
defparam fxp_functions_0_aadd_10_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a26.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_10_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_21_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a67.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_21_a67.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_19_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a62.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_19_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a21_sumout),
	.cout(fxp_functions_0_aadd_8_a22),
	.shareout());
defparam fxp_functions_0_aadd_8_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a21.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_8_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a57.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_17_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_6_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_15_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a52.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_15_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_6_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_6_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_6_a16_sumout),
	.cout(fxp_functions_0_aadd_6_a17),
	.shareout());
defparam fxp_functions_0_aadd_6_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_6_a16.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_6_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a47.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_13_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_4_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a_aq));
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_11_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a42.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_11_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_4_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_4_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_4_a11_sumout),
	.cout(fxp_functions_0_aadd_4_a12),
	.shareout());
defparam fxp_functions_0_aadd_4_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_4_a11.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_4_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a37.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_9_a37.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a32.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_7_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_5_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_5_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_5_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a27.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_5_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_3_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_3_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_3_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a22.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_3_a22.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_13_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_14_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_14_a41_sumout),
	.cout(fxp_functions_0_aadd_14_a42),
	.shareout());
defparam fxp_functions_0_aadd_14_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a41.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_14_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_15_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_16_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_16_a46_sumout),
	.cout(fxp_functions_0_aadd_16_a47),
	.shareout());
defparam fxp_functions_0_aadd_16_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a46.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_16_a46.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_17_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_18_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_18_a51_sumout),
	.cout(fxp_functions_0_aadd_18_a52),
	.shareout());
defparam fxp_functions_0_aadd_18_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a51.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_18_a51.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_19_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_20_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_20_a56_sumout),
	.cout(fxp_functions_0_aadd_20_a57),
	.shareout());
defparam fxp_functions_0_aadd_20_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a56.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_20_a56.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_21_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_22_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_22_a61_sumout),
	.cout(fxp_functions_0_aadd_22_a62),
	.shareout());
defparam fxp_functions_0_aadd_22_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a61.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_22_a61.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_23_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_24_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_24_a66_sumout),
	.cout(fxp_functions_0_aadd_24_a67),
	.shareout());
defparam fxp_functions_0_aadd_24_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a66.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_24_a66.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_25_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_26_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_26_a71_sumout),
	.cout(fxp_functions_0_aadd_26_a72),
	.shareout());
defparam fxp_functions_0_aadd_26_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a71.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_26_a71.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_27_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_28_a82_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_28_a76_sumout),
	.cout(fxp_functions_0_aadd_28_a77),
	.shareout());
defparam fxp_functions_0_aadd_28_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a76.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_28_a76.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a92(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_29_a92_cout),
	.shareout());
defparam fxp_functions_0_aadd_29_a92.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a92.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_29_a92.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_29_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_30_a87_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_30_a81_sumout),
	.cout(fxp_functions_0_aadd_30_a82),
	.shareout());
defparam fxp_functions_0_aadd_30_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a81.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_30_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_11_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a36_sumout),
	.cout(fxp_functions_0_aadd_12_a37),
	.shareout());
defparam fxp_functions_0_aadd_12_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a36.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a87(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_27_a87_cout),
	.shareout());
defparam fxp_functions_0_aadd_27_a87.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a87.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_27_a87.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a82(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_25_a82_cout),
	.shareout());
defparam fxp_functions_0_aadd_25_a82.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a82.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_25_a82.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_9_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_10_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_10_a31_sumout),
	.cout(fxp_functions_0_aadd_10_a32),
	.shareout());
defparam fxp_functions_0_aadd_10_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a31.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_10_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_23_a77_cout),
	.shareout());
defparam fxp_functions_0_aadd_23_a77.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a77.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_23_a77.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_21_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_21_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a72.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_21_a72.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_7_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a26_sumout),
	.cout(fxp_functions_0_aadd_8_a27),
	.shareout());
defparam fxp_functions_0_aadd_8_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a26.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_19_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_19_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a67.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_19_a67.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a62.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_17_a62.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_6_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(!fxp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_6_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_6_a21_sumout),
	.cout(fxp_functions_0_aadd_6_a22),
	.shareout());
defparam fxp_functions_0_aadd_6_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_6_a21.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_6_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_15_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_15_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a57.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_15_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a_aq));
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a52.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_13_a52.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_4_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a_aq),
	.datad(!fxp_functions_0_aadd_3_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_4_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_4_a16_sumout),
	.cout(fxp_functions_0_aadd_4_a17),
	.shareout());
defparam fxp_functions_0_aadd_4_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_4_a16.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_4_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_11_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_11_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a47.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_11_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a(
	.clk(clk),
	.d(radical[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a29_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a42.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_9_a42.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_7_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_7_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a37.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_7_a37.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_5_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_5_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a32.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_5_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_3_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_3_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a27.lut_mask = 64'h000000000F0FF0F0;
defparam fxp_functions_0_aadd_3_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_sM_opls_uid81_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_14_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_14_a47_cout),
	.shareout());
defparam fxp_functions_0_aadd_14_a47.extended_lut = "off";
defparam fxp_functions_0_aadd_14_a47.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_14_a47.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_sM_opls_uid91_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_16_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_16_a52_cout),
	.shareout());
defparam fxp_functions_0_aadd_16_a52.extended_lut = "off";
defparam fxp_functions_0_aadd_16_a52.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_16_a52.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_sM_opls_uid101_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_18_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_18_a57_cout),
	.shareout());
defparam fxp_functions_0_aadd_18_a57.extended_lut = "off";
defparam fxp_functions_0_aadd_18_a57.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_18_a57.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_sM_opls_uid111_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_20_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_20_a62_cout),
	.shareout());
defparam fxp_functions_0_aadd_20_a62.extended_lut = "off";
defparam fxp_functions_0_aadd_20_a62.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_20_a62.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_sM_opls_uid121_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_22_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_22_a67_cout),
	.shareout());
defparam fxp_functions_0_aadd_22_a67.extended_lut = "off";
defparam fxp_functions_0_aadd_22_a67.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_22_a67.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_sM_opls_uid131_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_24_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_24_a72_cout),
	.shareout());
defparam fxp_functions_0_aadd_24_a72.extended_lut = "off";
defparam fxp_functions_0_aadd_24_a72.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_24_a72.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_sM_opls_uid141_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_26_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_26_a77_cout),
	.shareout());
defparam fxp_functions_0_aadd_26_a77.extended_lut = "off";
defparam fxp_functions_0_aadd_26_a77.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_26_a77.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_sM_opls_uid151_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_28_a82(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_28_a82_cout),
	.shareout());
defparam fxp_functions_0_aadd_28_a82.extended_lut = "off";
defparam fxp_functions_0_aadd_28_a82.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_28_a82.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_sM_opls_uid161_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_30_a87(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_30_a87_cout),
	.shareout());
defparam fxp_functions_0_aadd_30_a87.extended_lut = "off";
defparam fxp_functions_0_aadd_30_a87.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_30_a87.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_sM_opls_uid71_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_12_a42_cout),
	.shareout());
defparam fxp_functions_0_aadd_12_a42.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a42.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_12_a42.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_sM_opls_uid61_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_10_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_10_a37_cout),
	.shareout());
defparam fxp_functions_0_aadd_10_a37.extended_lut = "off";
defparam fxp_functions_0_aadd_10_a37.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_10_a37.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_sM_opls_uid51_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_8_a32_cout),
	.shareout());
defparam fxp_functions_0_aadd_8_a32.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a32.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_8_a32.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a25_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a_aq));
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist25_sM_opls_uid41_sqrt_merged_bit_select_c_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_6_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_6_a27_cout),
	.shareout());
defparam fxp_functions_0_aadd_6_a27.extended_lut = "off";
defparam fxp_functions_0_aadd_6_a27.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_6_a27.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a27_a(
	.clk(clk),
	.d(radical[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a27_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a(
	.clk(clk),
	.d(radical[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a28_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_4_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_4_a22_cout),
	.shareout());
defparam fxp_functions_0_aadd_4_a22.extended_lut = "off";
defparam fxp_functions_0_aadd_4_a22.lut_mask = 64'h00000000FFFF0000;
defparam fxp_functions_0_aadd_4_a22.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_sM_opls_uid151_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a24_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a25_a(
	.clk(clk),
	.d(radical[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a25_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a26_a(
	.clk(clk),
	.d(radical[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a26_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_sM_opls_uid141_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a23_a(
	.clk(clk),
	.d(radical[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a24_a(
	.clk(clk),
	.d(radical[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a24_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_sM_opls_uid131_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a21_a(
	.clk(clk),
	.d(radical[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a22_a(
	.clk(clk),
	.d(radical[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(radical[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_sM_opls_uid121_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a20_a(
	.clk(clk),
	.d(radical[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(radical[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(radical[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_sM_opls_uid111_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(radical[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(radical[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_sM_opls_uid101_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(radical[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(radical[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_sM_opls_uid91_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(radical[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(radical[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(radical[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(radical[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_sM_opls_uid71_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(radical[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(radical[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_sM_opls_uid61_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(radical[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(radical[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_sM_opls_uid51_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(radical[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(radical[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist24_sM_opls_uid41_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(radical[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist26_sM_opls_uid21_sqrt_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aredist16_sM_opls_uid81_sqrt_merged_bit_select_b_1_q_a14_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_1_a0(
	.dataa(!radical[30]),
	.datab(!radical[28]),
	.datac(!radical[29]),
	.datad(!radical[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_1_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_1_a0.extended_lut = "off";
defparam fxp_functions_0_aadd_1_a0.lut_mask = 64'hD580D580D580D580;
defparam fxp_functions_0_aadd_1_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0(
	.dataa(!radical[30]),
	.datab(!radical[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_areduce_nor_0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_2_a0(
	.dataa(!fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq),
	.datab(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a0_a_aq),
	.datae(!fxp_functions_0_aredist27_sM_opls_uid21_sqrt_merged_bit_select_c_1_q_a2_a_aq),
	.dataf(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_2_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_2_a0.extended_lut = "off";
defparam fxp_functions_0_aadd_2_a0.lut_mask = 64'hDFFF200075558AAA;
defparam fxp_functions_0_aadd_2_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0(
	.dataa(!fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq),
	.datab(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_asM_decrms1_uid24_sqrt_sM_choosems_uid26_sqrt_merged_b1_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0(
	.dataa(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aadd_3_a1_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0.extended_lut = "off";
defparam fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0.lut_mask = 64'h4444444444444444;
defparam fxp_functions_0_asM_decrms1_uid34_sqrt_sM_choosems_uid36_sqrt_merged_b1_a3_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai240_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist44_sM_combine_uid20_sqrt_q_1_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai240_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai240_a0.extended_lut = "off";
defparam fxp_functions_0_ai240_a0.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_ai240_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a0(
	.dataa(!radical[30]),
	.datab(!radical[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_0_a0.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a0.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_aadd_0_a0.shared_arith = "off";

fourteennm_lcell_comb a_aGND(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(a_aGND_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam a_aGND.extended_lut = "off";
defparam a_aGND.lut_mask = 64'h0000000000000000;
defparam a_aGND.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_11_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_11_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_11_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_11_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_11_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_11_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_13_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_13_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_13_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_13_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_15_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_15_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_15_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_15_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_17_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_17_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_17_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_17_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_19_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_19_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_19_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_19_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_19_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_19_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_21_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_21_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_21_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_21_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_21_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_21_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_23_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_23_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_23_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_23_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_23_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_23_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_25_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_25_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_25_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_25_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_25_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_25_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_27_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_27_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_27_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_27_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_27_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_27_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_29_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_29_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_29_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_29_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_29_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_29_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_3_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_3_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_3_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_3_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_3_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_3_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_5_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_5_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_5_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_5_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_5_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_5_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_7_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_7_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_7_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_7_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a1_wirecell(
	.dataa(!fxp_functions_0_aadd_9_a1_sumout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_9_a1_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_9_a1_wirecell.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a1_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aadd_9_a1_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell(
	.dataa(!fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_asE_cmpge_uid23_sqrt_o_a5_a_a_wirecell.shared_arith = "off";

assign result[31] = a_aGND_acombout;

assign result[28] = a_aGND_acombout;

assign result[27] = a_aGND_acombout;

assign result[26] = a_aGND_acombout;

assign result[25] = a_aGND_acombout;

assign result[24] = a_aGND_acombout;

assign result[23] = a_aGND_acombout;

assign result[22] = a_aGND_acombout;

assign result[21] = a_aGND_acombout;

assign result[20] = a_aGND_acombout;

assign result[19] = a_aGND_acombout;

assign result[18] = a_aGND_acombout;

assign result[17] = a_aGND_acombout;

assign result[29] = a_aGND_acombout;

assign result[30] = a_aGND_acombout;

assign result[2] = fxp_functions_0_aadd_32_a11_sumout;

assign result[3] = fxp_functions_0_aadd_32_a16_sumout;

assign result[0] = fxp_functions_0_aadd_32_a1_sumout;

assign result[4] = fxp_functions_0_aadd_32_a21_sumout;

assign result[5] = fxp_functions_0_aadd_32_a26_sumout;

assign result[6] = fxp_functions_0_aadd_32_a31_sumout;

assign result[7] = fxp_functions_0_aadd_32_a36_sumout;

assign result[8] = fxp_functions_0_aadd_32_a41_sumout;

assign result[9] = fxp_functions_0_aadd_32_a46_sumout;

assign result[10] = fxp_functions_0_aadd_32_a51_sumout;

assign result[11] = fxp_functions_0_aadd_32_a56_sumout;

assign result[12] = fxp_functions_0_aadd_32_a61_sumout;

assign result[13] = fxp_functions_0_aadd_32_a66_sumout;

assign result[1] = fxp_functions_0_aadd_32_a6_sumout;

assign result[14] = fxp_functions_0_aadd_32_a71_sumout;

assign result[15] = fxp_functions_0_aadd_32_a76_sumout;

assign result[16] = fxp_functions_0_aadd_32_a81_sumout;

endmodule
