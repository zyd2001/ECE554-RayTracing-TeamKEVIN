// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/20/2021 23:10:26"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Float_Div (
	q,
	clk,
	areset,
	en,
	b,
	a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	clk;
input 	areset;
input 	[0:0] en;
input 	[31:0] b;
input 	[31:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a0_a_aq;
wire fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist19_excI_x_uid27_fpDivTest_q_1_q_a0_a_aq;
wire fp_functions_0_aexpOvf_uid84_fpDivTest_o_a12_a_aq;
wire fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a_aq;
wire fp_functions_0_aredist17_excZ_y_uid37_fpDivTest_q_25_q_a0_a_aq;
wire fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist23_excZ_x_uid23_fpDivTest_q_25_q_a0_a_aq;
wire fp_functions_0_aexpUdf_uid81_fpDivTest_o_a12_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a8_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a9_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a10_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a11_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a12_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a13_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a14_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a15_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a16_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a17_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a18_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a19_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a20_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a21_a_aq;
wire fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a22_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aadd_16_a1_sumout;
wire fp_functions_0_aadd_16_a2;
wire fp_functions_0_aadd_17_a1_sumout;
wire fp_functions_0_aadd_18_a1_sumout;
wire fp_functions_0_aadd_16_a6_sumout;
wire fp_functions_0_aadd_16_a7;
wire fp_functions_0_aadd_16_a11_sumout;
wire fp_functions_0_aadd_16_a12;
wire fp_functions_0_aadd_16_a16_sumout;
wire fp_functions_0_aadd_16_a17;
wire fp_functions_0_aadd_16_a21_sumout;
wire fp_functions_0_aadd_16_a22;
wire fp_functions_0_aadd_16_a26_sumout;
wire fp_functions_0_aadd_16_a27;
wire fp_functions_0_aadd_16_a31_sumout;
wire fp_functions_0_aadd_16_a32;
wire fp_functions_0_aadd_16_a36_sumout;
wire fp_functions_0_aadd_16_a37;
wire fp_functions_0_aadd_16_a41_sumout;
wire fp_functions_0_aadd_16_a42;
wire fp_functions_0_aadd_16_a46_sumout;
wire fp_functions_0_aadd_16_a47;
wire fp_functions_0_aadd_16_a51_sumout;
wire fp_functions_0_aadd_16_a52;
wire fp_functions_0_aadd_16_a56_sumout;
wire fp_functions_0_aadd_16_a57;
wire fp_functions_0_aadd_16_a61_sumout;
wire fp_functions_0_aadd_16_a62;
wire fp_functions_0_aadd_16_a66_sumout;
wire fp_functions_0_aadd_16_a67;
wire fp_functions_0_aadd_16_a71_sumout;
wire fp_functions_0_aadd_16_a72;
wire fp_functions_0_aadd_16_a76_sumout;
wire fp_functions_0_aadd_16_a77;
wire fp_functions_0_aadd_16_a81_sumout;
wire fp_functions_0_aadd_16_a82;
wire fp_functions_0_aadd_16_a86_sumout;
wire fp_functions_0_aadd_16_a87;
wire fp_functions_0_aadd_16_a91_sumout;
wire fp_functions_0_aadd_16_a92;
wire fp_functions_0_aadd_16_a96_sumout;
wire fp_functions_0_aadd_16_a97;
wire fp_functions_0_aadd_16_a101_sumout;
wire fp_functions_0_aadd_16_a102;
wire fp_functions_0_aadd_16_a106_sumout;
wire fp_functions_0_aadd_16_a107;
wire fp_functions_0_aadd_16_a111_sumout;
wire fp_functions_0_aadd_16_a112;
wire fp_functions_0_aadd_16_a116_sumout;
wire fp_functions_0_aadd_16_a117;
wire fp_functions_0_aadd_16_a121_sumout;
wire fp_functions_0_aadd_16_a122;
wire fp_functions_0_aadd_16_a126_sumout;
wire fp_functions_0_aadd_16_a127;
wire fp_functions_0_aadd_16_a131_sumout;
wire fp_functions_0_aadd_16_a132;
wire fp_functions_0_aadd_16_a136_sumout;
wire fp_functions_0_aadd_16_a137;
wire fp_functions_0_aadd_16_a141_sumout;
wire fp_functions_0_aadd_16_a142;
wire fp_functions_0_aadd_16_a146_sumout;
wire fp_functions_0_aadd_16_a147;
wire fp_functions_0_aadd_16_a151_sumout;
wire fp_functions_0_aadd_16_a152;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a0_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a1_a_aq;
wire fp_functions_0_aadd_16_a156_sumout;
wire fp_functions_0_aadd_17_a7_cout;
wire fp_functions_0_aadd_18_a7_cout;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a2_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a3_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a4_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a5_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a6_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a7_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a8_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a9_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a10_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a11_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a12_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a13_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a14_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a15_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a16_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a17_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a18_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a19_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a20_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a21_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a22_a_aq;
wire fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a23_a_aq;
wire fp_functions_0_aredist5_norm_uid67_fpDivTest_b_1_q_a0_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a0_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a1_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a2_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a3_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a4_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a5_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a6_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a7_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a_aq;
wire fp_functions_0_aadd_16_a161_sumout;
wire fp_functions_0_aadd_16_a162;
wire fp_functions_0_aadd_17_a12_cout;
wire fp_functions_0_aadd_18_a12_cout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aadd_15_a1_sumout;
wire fp_functions_0_aadd_15_a2;
wire fp_functions_0_aadd_15_a6_sumout;
wire fp_functions_0_aadd_15_a7;
wire fp_functions_0_aadd_15_a11_sumout;
wire fp_functions_0_aadd_15_a12;
wire fp_functions_0_aadd_15_a16_sumout;
wire fp_functions_0_aadd_15_a17;
wire fp_functions_0_aadd_15_a21_sumout;
wire fp_functions_0_aadd_15_a22;
wire fp_functions_0_aadd_15_a26_sumout;
wire fp_functions_0_aadd_15_a27;
wire fp_functions_0_aadd_15_a31_sumout;
wire fp_functions_0_aadd_15_a32;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a24_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a25_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a26_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a27_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a28_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a29_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a30_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a31_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a32_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a33_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a34_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a35_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a36_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a37_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a38_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a39_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a40_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a41_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a42_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a43_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a44_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a45_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a46_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a47_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a48_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a49_a;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a23_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aadd_15_a36_sumout;
wire fp_functions_0_aadd_16_a166_sumout;
wire fp_functions_0_aadd_16_a167;
wire fp_functions_0_aadd_17_a17_cout;
wire fp_functions_0_aadd_18_a17_cout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aadd_15_a41_sumout;
wire fp_functions_0_aadd_15_a42;
wire fp_functions_0_aexpR_uid48_fpDivTest_o_a8_a_aq;
wire fp_functions_0_aadd_17_a22_cout;
wire fp_functions_0_aadd_18_a22_cout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a0_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a1_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a2_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a3_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a4_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a5_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a6_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a7_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a8_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a9_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a10_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a11_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a12_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a13_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a14_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a15_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a16_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a17_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a18_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a19_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a20_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a21_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a22_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a23_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a24_a_aq;
wire fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a25_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aadd_17_a27_cout;
wire fp_functions_0_aadd_18_a27_cout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_afracXIsZero_uid25_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq;
wire fp_functions_0_aadd_11_a1_sumout;
wire fp_functions_0_aadd_11_a2;
wire fp_functions_0_aadd_11_a6_sumout;
wire fp_functions_0_aadd_11_a7;
wire fp_functions_0_aadd_11_a11_sumout;
wire fp_functions_0_aadd_11_a12;
wire fp_functions_0_aadd_11_a16_sumout;
wire fp_functions_0_aadd_11_a17;
wire fp_functions_0_aadd_11_a21_sumout;
wire fp_functions_0_aadd_11_a22;
wire fp_functions_0_aadd_11_a26_sumout;
wire fp_functions_0_aadd_11_a27;
wire fp_functions_0_aadd_11_a31_sumout;
wire fp_functions_0_aadd_11_a32;
wire fp_functions_0_aadd_11_a36_sumout;
wire fp_functions_0_aadd_11_a37;
wire fp_functions_0_aadd_11_a41_sumout;
wire fp_functions_0_aadd_11_a42;
wire fp_functions_0_aadd_11_a46_sumout;
wire fp_functions_0_aadd_11_a47;
wire fp_functions_0_aadd_11_a51_sumout;
wire fp_functions_0_aadd_11_a52;
wire fp_functions_0_aadd_11_a56_sumout;
wire fp_functions_0_aadd_11_a57;
wire fp_functions_0_aadd_11_a61_sumout;
wire fp_functions_0_aadd_11_a62;
wire fp_functions_0_aadd_11_a66_sumout;
wire fp_functions_0_aadd_11_a67;
wire fp_functions_0_aadd_11_a71_sumout;
wire fp_functions_0_aadd_11_a72;
wire fp_functions_0_aadd_11_a76_sumout;
wire fp_functions_0_aadd_11_a77;
wire fp_functions_0_aadd_11_a81_sumout;
wire fp_functions_0_aadd_11_a82;
wire fp_functions_0_aadd_11_a86_sumout;
wire fp_functions_0_aadd_11_a87;
wire fp_functions_0_aadd_11_a91_sumout;
wire fp_functions_0_aadd_11_a92;
wire fp_functions_0_aadd_11_a96_sumout;
wire fp_functions_0_aadd_11_a97;
wire fp_functions_0_aadd_11_a101_sumout;
wire fp_functions_0_aadd_11_a102;
wire fp_functions_0_aadd_11_a106_sumout;
wire fp_functions_0_aadd_11_a107;
wire fp_functions_0_aadd_11_a111_sumout;
wire fp_functions_0_aadd_11_a112;
wire fp_functions_0_aadd_11_a116_sumout;
wire fp_functions_0_aadd_11_a117;
wire fp_functions_0_aadd_11_a121_sumout;
wire fp_functions_0_aadd_11_a122;
wire fp_functions_0_aadd_11_a126_sumout;
wire fp_functions_0_aadd_11_a127;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq_aq;
wire fp_functions_0_aadd_17_a32_cout;
wire fp_functions_0_aadd_18_a32_cout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq_aq;
wire fp_functions_0_aadd_14_a1_sumout;
wire fp_functions_0_aadd_14_a2;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a1_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a2_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a3_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a4_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a5_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a6_a_aq;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a7_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_aadd_11_a132_cout;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a;
wire fp_functions_0_aexpXmY_uid47_fpDivTest_o_a8_a_aq;
wire fp_functions_0_aadd_17_a37_cout;
wire fp_functions_0_aadd_18_a37_cout;
wire fp_functions_0_aadd_14_a7_cout;
wire fp_functions_0_aadd_14_a11_sumout;
wire fp_functions_0_aadd_14_a12;
wire fp_functions_0_aadd_14_a16_sumout;
wire fp_functions_0_aadd_14_a17;
wire fp_functions_0_aadd_14_a21_sumout;
wire fp_functions_0_aadd_14_a22;
wire fp_functions_0_aadd_14_a26_sumout;
wire fp_functions_0_aadd_14_a27;
wire fp_functions_0_aadd_14_a31_sumout;
wire fp_functions_0_aadd_14_a32;
wire fp_functions_0_aadd_14_a36_sumout;
wire fp_functions_0_aadd_14_a37;
wire fp_functions_0_aadd_14_a41_sumout;
wire fp_functions_0_aadd_14_a42;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_afracYPostZ_uid56_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmpReg_q_a0_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a24_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a25_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a26_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a27_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a28_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a29_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a30_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a31_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a32_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a33_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a34_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a35_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a36_a;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_aadd_11_a137_cout;
wire fp_functions_0_aadd_14_a46_sumout;
wire fp_functions_0_aadd_17_a42_cout;
wire fp_functions_0_aadd_18_a42_cout;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aadd_11_a141_sumout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_aadd_11_a147_cout;
wire fp_functions_0_aadd_17_a47_cout;
wire fp_functions_0_aadd_18_a47_cout;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a29_a;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq_aq;
wire fp_functions_0_aredist2_lowRangeB_uid126_invPolyEval_b_1_q_a0_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a0_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a1_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a2_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a3_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a4_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a5_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a6_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a7_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a8_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a9_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a10_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a11_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a12_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a13_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a14_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a15_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a16_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a17_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a18_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a19_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a20_a_aq;
wire fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a21_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a8_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a9_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a10_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a11_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a12_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a13_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_aadd_17_a52_cout;
wire fp_functions_0_aadd_18_a52_cout;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aadd_6_a1_sumout;
wire fp_functions_0_aadd_6_a2;
wire fp_functions_0_aadd_6_a6_sumout;
wire fp_functions_0_aadd_6_a7;
wire fp_functions_0_aadd_6_a11_sumout;
wire fp_functions_0_aadd_6_a12;
wire fp_functions_0_aadd_6_a16_sumout;
wire fp_functions_0_aadd_6_a17;
wire fp_functions_0_aadd_6_a21_sumout;
wire fp_functions_0_aadd_6_a22;
wire fp_functions_0_aadd_6_a26_sumout;
wire fp_functions_0_aadd_6_a27;
wire fp_functions_0_aadd_6_a31_sumout;
wire fp_functions_0_aadd_6_a32;
wire fp_functions_0_aadd_6_a36_sumout;
wire fp_functions_0_aadd_6_a37;
wire fp_functions_0_aadd_6_a41_sumout;
wire fp_functions_0_aadd_6_a42;
wire fp_functions_0_aadd_6_a46_sumout;
wire fp_functions_0_aadd_6_a47;
wire fp_functions_0_aadd_6_a51_sumout;
wire fp_functions_0_aadd_6_a52;
wire fp_functions_0_aadd_6_a56_sumout;
wire fp_functions_0_aadd_6_a57;
wire fp_functions_0_aadd_6_a61_sumout;
wire fp_functions_0_aadd_6_a62;
wire fp_functions_0_aadd_6_a66_sumout;
wire fp_functions_0_aadd_6_a67;
wire fp_functions_0_aadd_6_a71_sumout;
wire fp_functions_0_aadd_6_a72;
wire fp_functions_0_aadd_6_a76_sumout;
wire fp_functions_0_aadd_6_a77;
wire fp_functions_0_aadd_6_a81_sumout;
wire fp_functions_0_aadd_6_a82;
wire fp_functions_0_aadd_6_a86_sumout;
wire fp_functions_0_aadd_6_a87;
wire fp_functions_0_aadd_6_a91_sumout;
wire fp_functions_0_aadd_6_a92;
wire fp_functions_0_aadd_6_a96_sumout;
wire fp_functions_0_aadd_6_a97;
wire fp_functions_0_aadd_6_a101_sumout;
wire fp_functions_0_aadd_6_a102;
wire fp_functions_0_aadd_6_a106_sumout;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA24;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA25;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA26;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA27;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA28;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA29;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA30;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA31;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA32;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA33;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA34;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA35;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA36;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a0_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a1_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a2_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a3_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a4_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a5_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a6_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a7_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a8_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a9_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a10_a_aq;
wire fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a11_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a0_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a2_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a3_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a4_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a5_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a6_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a7_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a8_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a9_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a10_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a11_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a12_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a13_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a0_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_cmpReg_q_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a16_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a2_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a3_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a4_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a5_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a6_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a7_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a8_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a9_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a10_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a11_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a12_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a13_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a0_a_aq;
wire fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a17_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a18_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a19_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a20_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a21_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a22_a_a0_a_aq;
wire fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq;
wire fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq;
wire fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a23_a_a0_a_aq;
wire fp_functions_0_aexcZ_x_uid23_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aexcZ_y_uid37_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aexpXIsMax_uid38_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_afracXIsZero_uid39_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aexpXIsMax_uid24_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_asignR_uid46_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_afracYZero_uid15_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout;
wire fp_functions_0_aMux_31_a0_combout;
wire fp_functions_0_aMux_32_a2_combout;
wire fp_functions_0_aMux_31_a1_combout;
wire fp_functions_0_aMux_30_a0_combout;
wire fp_functions_0_aMux_29_a0_combout;
wire fp_functions_0_aMux_28_a0_combout;
wire fp_functions_0_aMux_27_a0_combout;
wire fp_functions_0_aMux_26_a0_combout;
wire fp_functions_0_aMux_25_a0_combout;
wire fp_functions_0_aMux_24_a0_combout;
wire fp_functions_0_aMux_23_a0_combout;
wire fp_functions_0_aMux_22_a0_combout;
wire fp_functions_0_aMux_21_a0_combout;
wire fp_functions_0_aMux_20_a0_combout;
wire fp_functions_0_aMux_19_a0_combout;
wire fp_functions_0_aMux_18_a0_combout;
wire fp_functions_0_aMux_17_a0_combout;
wire fp_functions_0_aMux_16_a0_combout;
wire fp_functions_0_aMux_15_a0_combout;
wire fp_functions_0_aMux_14_a0_combout;
wire fp_functions_0_aMux_13_a0_combout;
wire fp_functions_0_aMux_12_a0_combout;
wire fp_functions_0_aMux_11_a0_combout;
wire fp_functions_0_aMux_10_a0_combout;
wire fp_functions_0_aMux_9_a2_combout;
wire fp_functions_0_aMux_9_a3_combout;
wire fp_functions_0_aMux_9_a4_combout;
wire fp_functions_0_aMux_9_a5_combout;
wire fp_functions_0_aMux_9_a6_combout;
wire fp_functions_0_aMux_9_a7_combout;
wire fp_functions_0_aMux_9_a8_combout;
wire fp_functions_0_aMux_9_a9_combout;
wire fp_functions_0_adivR_uid110_fpDivTest_q_a31_a_acombout;
wire fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1_combout;
wire fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout;
wire fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a_acombout;
wire fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a_acombout;
wire fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a_acombout;
wire fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fp_functions_0_ai2642_a0_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fp_functions_0_ai2642_a1_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout;
wire fp_functions_0_ai2690_a0_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fp_functions_0_ai2690_a1_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fp_functions_0_ai2690_a2_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fp_functions_0_ai2690_a3_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fp_functions_0_ai2690_a4_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fp_functions_0_ai2690_a5_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fp_functions_0_ai2690_a6_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fp_functions_0_ai2690_a7_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fp_functions_0_ai2690_a8_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a_aq;
wire fp_functions_0_ai2690_a9_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a_aq;
wire fp_functions_0_ai2690_a10_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a_aq;
wire fp_functions_0_ai2690_a11_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a_aq;
wire fp_functions_0_ai2690_a12_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a_aq;
wire fp_functions_0_ai2690_a13_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a_aq;
wire fp_functions_0_ai2690_a14_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a_aq;
wire fp_functions_0_ai2690_a15_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a_aq;
wire fp_functions_0_ai2690_a16_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a_aq;
wire fp_functions_0_ai2690_a17_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a_aq;
wire fp_functions_0_ai2690_a18_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a_aq;
wire fp_functions_0_ai2690_a19_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a_aq;
wire fp_functions_0_ai2690_a20_combout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a48_a_aq;
wire fp_functions_0_ai2690_a21_combout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a23_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a23_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a24_a_aq;
wire fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a25_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai401_a0_combout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq;
wire fp_functions_0_ai2307_a0_combout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai456_a0_combout;
wire fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_8_acombout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0_combout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1_combout;
wire fp_functions_0_ai2418_a0_combout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2_combout;
wire fp_functions_0_ai2418_a1_combout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3_combout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4_combout;
wire fp_functions_0_areduce_nor_20_acombout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_ai413_a0_combout;
wire fp_functions_0_ai413_a1_combout;
wire fp_functions_0_ai413_a2_combout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_ai2329_a0_combout;
wire fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0_combout;
wire fp_functions_0_aadd_13_a0_combout;
wire fp_functions_0_ai2329_a1_combout;
wire fp_functions_0_ai2329_a2_combout;
wire fp_functions_0_ai2329_a3_combout;
wire fp_functions_0_areduce_nor_4_a0_combout;
wire fp_functions_0_areduce_nor_4_a1_combout;
wire fp_functions_0_areduce_nor_4_a2_combout;
wire fp_functions_0_areduce_nor_4_acombout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq;
wire fp_functions_0_areduce_nor_9_acombout;
wire fp_functions_0_areduce_nor_18_acombout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq;
wire fp_functions_0_ai119_a0_combout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a_acombout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0_combout;
wire fp_functions_0_ai182_a0_combout;
wire fp_functions_0_ai182_a1_combout;
wire fp_functions_0_ai182_a2_combout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1_combout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2_combout;
wire fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3_combout;
wire fp_functions_0_areduce_nor_19_acombout;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fp_functions_0_ai134_a0_combout;
wire fp_functions_0_ai138_a0_combout;
wire fp_functions_0_ai138_a1_combout;
wire fp_functions_0_ai138_a2_combout;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fp_functions_0_areduce_nor_3_acombout;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai1513_a0_combout;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai1544_a0_combout;
wire fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_14_acombout;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai1191_a0_combout;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fp_functions_0_ai1525_a0_combout;
wire fp_functions_0_ai1525_a1_combout;
wire fp_functions_0_ai1525_a2_combout;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai1222_a0_combout;
wire fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_12_acombout;
wire fp_functions_0_areduce_nor_15_acombout;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout;
wire fp_functions_0_ai1203_a0_combout;
wire fp_functions_0_ai1203_a1_combout;
wire fp_functions_0_ai1203_a2_combout;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_ai899_a0_combout;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_areduce_nor_13_acombout;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0_combout;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1_combout;
wire fp_functions_0_ai930_a0_combout;
wire fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2_combout;
wire fp_functions_0_areduce_nor_10_acombout;
wire fp_functions_0_ai911_a0_combout;
wire fp_functions_0_ai911_a1_combout;
wire fp_functions_0_ai911_a2_combout;
wire fp_functions_0_areduce_nor_11_acombout;
wire fp_functions_0_areduce_nor_7_a0_combout;
wire fp_functions_0_areduce_nor_7_acombout;
wire fp_functions_0_areduce_nor_6_a0_combout;
wire fp_functions_0_areduce_nor_6_acombout;
wire fp_functions_0_areduce_nor_1_a0_combout;
wire fp_functions_0_areduce_nor_1_acombout;
wire fp_functions_0_areduce_nor_16_a0_combout;
wire fp_functions_0_areduce_nor_16_a1_combout;
wire fp_functions_0_areduce_nor_16_a2_combout;
wire fp_functions_0_areduce_nor_16_a3_combout;
wire fp_functions_0_areduce_nor_16_acombout;
wire fp_functions_0_areduce_nor_5_a0_combout;
wire fp_functions_0_areduce_nor_5_acombout;
wire fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a_acombout;
wire fp_functions_0_areduce_nor_4_a3_combout;
wire fp_functions_0_areduce_nor_4_a4_combout;

wire [63:0] fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus;
wire [63:0] fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [63:0] fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;

assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a0_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a1_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a2_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a3_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a4_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a5_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a6_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a7_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a8_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a9_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a10_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a11_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a12_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a13_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a14_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a15_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a16_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a17_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a18_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a19_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a20_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a21_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a22_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a23_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a24_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a25_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a26_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a27_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a28_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a29_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a30_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a31_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a32_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a33_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a34_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a35_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a36_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a37_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a38_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a39_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a40_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a41_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a42_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a43_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a44_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a45_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a46_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a47_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a48_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a49_a = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a23_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19 = fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19 = fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus[0];

assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a0_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a1_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a2_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a3_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a4_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a5_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a6_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a7_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a8_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a9_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a10_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a11_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a12_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a13_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a14_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a15_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a16_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a17_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a18_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a19_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a20_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a21_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a22_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a23_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a24_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a25_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a26_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a27_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a28_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a29_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a30_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a31_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a32_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a33_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a34_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a35_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a36_a = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA37 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA38 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA39 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA40 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA41 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA42 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA43 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA44 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA45 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA46 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA47 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA48 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA49 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a29_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a0_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a1_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a2_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a3_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a4_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a5_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a6_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a7_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a8_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a9_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a10_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a11_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a12_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a13_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a14_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a15_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a16_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a17_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a18_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a19_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a20_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a21_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a22_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a23_a = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA24 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA25 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA26 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA27 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA28 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA29 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA30 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA31 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA32 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA33 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA34 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA35 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA36 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA37 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA38 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA39 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA40 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA41 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA42 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA43 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA44 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA45 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA46 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA47 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA48 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA49 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

fourteennm_ff fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist19_excI_x_uid27_fpDivTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist19_excI_x_uid27_fpDivTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist19_excI_x_uid27_fpDivTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist19_excI_x_uid27_fpDivTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpOvf_uid84_fpDivTest_o_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_17_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpOvf_uid84_fpDivTest_o_a12_a_aq));
defparam fp_functions_0_aexpOvf_uid84_fpDivTest_o_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpOvf_uid84_fpDivTest_o_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_excZ_y_uid37_fpDivTest_q_25_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_excZ_y_uid37_fpDivTest_q_25_q_a0_a_aq));
defparam fp_functions_0_aredist17_excZ_y_uid37_fpDivTest_q_25_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_excZ_y_uid37_fpDivTest_q_25_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist23_excZ_x_uid23_fpDivTest_q_25_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist23_excZ_x_uid23_fpDivTest_q_25_q_a0_a_aq));
defparam fp_functions_0_aredist23_excZ_x_uid23_fpDivTest_q_25_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist23_excZ_x_uid23_fpDivTest_q_25_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpUdf_uid81_fpDivTest_o_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_18_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpUdf_uid81_fpDivTest_o_a12_a_aq));
defparam fp_functions_0_aexpUdf_uid81_fpDivTest_o_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpUdf_uid81_fpDivTest_o_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_16_a151_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_16_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a0_a_aq),
	.datad(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a1_sumout),
	.cout(fp_functions_0_aadd_16_a2),
	.shareout());
defparam fp_functions_0_aadd_16_a1.extended_lut = "off";
defparam fp_functions_0_aadd_16_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_16_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_17_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a156_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_17_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_17_a1.extended_lut = "off";
defparam fp_functions_0_aadd_17_a1.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_17_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a156_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_18_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_18_a1.extended_lut = "off";
defparam fp_functions_0_aadd_18_a1.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a6_sumout),
	.cout(fp_functions_0_aadd_16_a7),
	.shareout());
defparam fp_functions_0_aadd_16_a6.extended_lut = "off";
defparam fp_functions_0_aadd_16_a6.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a11_sumout),
	.cout(fp_functions_0_aadd_16_a12),
	.shareout());
defparam fp_functions_0_aadd_16_a11.extended_lut = "off";
defparam fp_functions_0_aadd_16_a11.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a16_sumout),
	.cout(fp_functions_0_aadd_16_a17),
	.shareout());
defparam fp_functions_0_aadd_16_a16.extended_lut = "off";
defparam fp_functions_0_aadd_16_a16.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a21_sumout),
	.cout(fp_functions_0_aadd_16_a22),
	.shareout());
defparam fp_functions_0_aadd_16_a21.extended_lut = "off";
defparam fp_functions_0_aadd_16_a21.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a26_sumout),
	.cout(fp_functions_0_aadd_16_a27),
	.shareout());
defparam fp_functions_0_aadd_16_a26.extended_lut = "off";
defparam fp_functions_0_aadd_16_a26.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a31_sumout),
	.cout(fp_functions_0_aadd_16_a32),
	.shareout());
defparam fp_functions_0_aadd_16_a31.extended_lut = "off";
defparam fp_functions_0_aadd_16_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a36_sumout),
	.cout(fp_functions_0_aadd_16_a37),
	.shareout());
defparam fp_functions_0_aadd_16_a36.extended_lut = "off";
defparam fp_functions_0_aadd_16_a36.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a41_sumout),
	.cout(fp_functions_0_aadd_16_a42),
	.shareout());
defparam fp_functions_0_aadd_16_a41.extended_lut = "off";
defparam fp_functions_0_aadd_16_a41.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a46_sumout),
	.cout(fp_functions_0_aadd_16_a47),
	.shareout());
defparam fp_functions_0_aadd_16_a46.extended_lut = "off";
defparam fp_functions_0_aadd_16_a46.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a51_sumout),
	.cout(fp_functions_0_aadd_16_a52),
	.shareout());
defparam fp_functions_0_aadd_16_a51.extended_lut = "off";
defparam fp_functions_0_aadd_16_a51.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a56_sumout),
	.cout(fp_functions_0_aadd_16_a57),
	.shareout());
defparam fp_functions_0_aadd_16_a56.extended_lut = "off";
defparam fp_functions_0_aadd_16_a56.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a61_sumout),
	.cout(fp_functions_0_aadd_16_a62),
	.shareout());
defparam fp_functions_0_aadd_16_a61.extended_lut = "off";
defparam fp_functions_0_aadd_16_a61.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a66_sumout),
	.cout(fp_functions_0_aadd_16_a67),
	.shareout());
defparam fp_functions_0_aadd_16_a66.extended_lut = "off";
defparam fp_functions_0_aadd_16_a66.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a71_sumout),
	.cout(fp_functions_0_aadd_16_a72),
	.shareout());
defparam fp_functions_0_aadd_16_a71.extended_lut = "off";
defparam fp_functions_0_aadd_16_a71.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a76_sumout),
	.cout(fp_functions_0_aadd_16_a77),
	.shareout());
defparam fp_functions_0_aadd_16_a76.extended_lut = "off";
defparam fp_functions_0_aadd_16_a76.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a81_sumout),
	.cout(fp_functions_0_aadd_16_a82),
	.shareout());
defparam fp_functions_0_aadd_16_a81.extended_lut = "off";
defparam fp_functions_0_aadd_16_a81.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a86_sumout),
	.cout(fp_functions_0_aadd_16_a87),
	.shareout());
defparam fp_functions_0_aadd_16_a86.extended_lut = "off";
defparam fp_functions_0_aadd_16_a86.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a91_sumout),
	.cout(fp_functions_0_aadd_16_a92),
	.shareout());
defparam fp_functions_0_aadd_16_a91.extended_lut = "off";
defparam fp_functions_0_aadd_16_a91.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a96_sumout),
	.cout(fp_functions_0_aadd_16_a97),
	.shareout());
defparam fp_functions_0_aadd_16_a96.extended_lut = "off";
defparam fp_functions_0_aadd_16_a96.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a101_sumout),
	.cout(fp_functions_0_aadd_16_a102),
	.shareout());
defparam fp_functions_0_aadd_16_a101.extended_lut = "off";
defparam fp_functions_0_aadd_16_a101.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a106_sumout),
	.cout(fp_functions_0_aadd_16_a107),
	.shareout());
defparam fp_functions_0_aadd_16_a106.extended_lut = "off";
defparam fp_functions_0_aadd_16_a106.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a111_sumout),
	.cout(fp_functions_0_aadd_16_a112),
	.shareout());
defparam fp_functions_0_aadd_16_a111.extended_lut = "off";
defparam fp_functions_0_aadd_16_a111.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist5_norm_uid67_fpDivTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aexpR_uid48_fpDivTest_o_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a116_sumout),
	.cout(fp_functions_0_aadd_16_a117),
	.shareout());
defparam fp_functions_0_aadd_16_a116.extended_lut = "off";
defparam fp_functions_0_aadd_16_a116.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_16_a116.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a121_sumout),
	.cout(fp_functions_0_aadd_16_a122),
	.shareout());
defparam fp_functions_0_aadd_16_a121.extended_lut = "off";
defparam fp_functions_0_aadd_16_a121.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a121.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a126_sumout),
	.cout(fp_functions_0_aadd_16_a127),
	.shareout());
defparam fp_functions_0_aadd_16_a126.extended_lut = "off";
defparam fp_functions_0_aadd_16_a126.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a126.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a131_sumout),
	.cout(fp_functions_0_aadd_16_a132),
	.shareout());
defparam fp_functions_0_aadd_16_a131.extended_lut = "off";
defparam fp_functions_0_aadd_16_a131.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a131.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a136_sumout),
	.cout(fp_functions_0_aadd_16_a137),
	.shareout());
defparam fp_functions_0_aadd_16_a136.extended_lut = "off";
defparam fp_functions_0_aadd_16_a136.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a136.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a141_sumout),
	.cout(fp_functions_0_aadd_16_a142),
	.shareout());
defparam fp_functions_0_aadd_16_a141.extended_lut = "off";
defparam fp_functions_0_aadd_16_a141.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a141.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a146_sumout),
	.cout(fp_functions_0_aadd_16_a147),
	.shareout());
defparam fp_functions_0_aadd_16_a146.extended_lut = "off";
defparam fp_functions_0_aadd_16_a146.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a146.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a151_sumout),
	.cout(fp_functions_0_aadd_16_a152),
	.shareout());
defparam fp_functions_0_aadd_16_a151.extended_lut = "off";
defparam fp_functions_0_aadd_16_a151.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a151.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai2642_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a0_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai2642_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a1_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_16_a156(
	.dataa(!fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a162),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a156_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_16_a156.extended_lut = "off";
defparam fp_functions_0_aadd_16_a156.lut_mask = 64'h0000000000005555;
defparam fp_functions_0_aadd_16_a156.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_17_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a156_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a7.extended_lut = "off";
defparam fp_functions_0_aadd_17_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_17_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a156_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a7.extended_lut = "off";
defparam fp_functions_0_aadd_18_a7.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a7.shared_arith = "off";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a2_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a3_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a4_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a5_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a6_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a7_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a8_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a9_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a10_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a11_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a12_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a13_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a14_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a15_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a16_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a17_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a18_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a17_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a19_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a18_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a20_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a19_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a21_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a20_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a22_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai2690_a21_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a23_a_aq));
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_anormFracRnd_uid70_fpDivTest_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_norm_uid67_fpDivTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_norm_uid67_fpDivTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist5_norm_uid67_fpDivTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_norm_uid67_fpDivTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a0_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a1_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a2_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a3_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a4_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a5_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a6_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a7_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_16_a161(
	.dataa(!fp_functions_0_aexpR_uid48_fpDivTest_o_a9_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a167),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a161_sumout),
	.cout(fp_functions_0_aadd_16_a162),
	.shareout());
defparam fp_functions_0_aadd_16_a161.extended_lut = "off";
defparam fp_functions_0_aadd_16_a161.lut_mask = 64'h0000000000005555;
defparam fp_functions_0_aadd_16_a161.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_17_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a161_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a12.extended_lut = "off";
defparam fp_functions_0_aadd_17_a12.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_17_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a161_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a12.extended_lut = "off";
defparam fp_functions_0_aadd_18_a12.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a12.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_15_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a1_sumout),
	.cout(fp_functions_0_aadd_15_a2),
	.shareout());
defparam fp_functions_0_aadd_15_a1.extended_lut = "off";
defparam fp_functions_0_aadd_15_a1.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_15_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_15_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a6_sumout),
	.cout(fp_functions_0_aadd_15_a7),
	.shareout());
defparam fp_functions_0_aadd_15_a6.extended_lut = "off";
defparam fp_functions_0_aadd_15_a6.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_15_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_15_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a11_sumout),
	.cout(fp_functions_0_aadd_15_a12),
	.shareout());
defparam fp_functions_0_aadd_15_a11.extended_lut = "off";
defparam fp_functions_0_aadd_15_a11.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_15_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_15_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a16_sumout),
	.cout(fp_functions_0_aadd_15_a17),
	.shareout());
defparam fp_functions_0_aadd_15_a16.extended_lut = "off";
defparam fp_functions_0_aadd_15_a16.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_15_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_15_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a21_sumout),
	.cout(fp_functions_0_aadd_15_a22),
	.shareout());
defparam fp_functions_0_aadd_15_a21.extended_lut = "off";
defparam fp_functions_0_aadd_15_a21.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_15_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_15_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a26_sumout),
	.cout(fp_functions_0_aadd_15_a27),
	.shareout());
defparam fp_functions_0_aadd_15_a26.extended_lut = "off";
defparam fp_functions_0_aadd_15_a26.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_15_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_15_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a31_sumout),
	.cout(fp_functions_0_aadd_15_a32),
	.shareout());
defparam fp_functions_0_aadd_15_a31.extended_lut = "off";
defparam fp_functions_0_aadd_15_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_15_a31.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a23_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a22_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a21_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a20_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a19_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a18_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a17_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a16_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a15_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a14_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a13_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a12_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a25_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a24_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a23_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a22_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a21_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a20_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a19_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a18_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a17_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a16_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a15_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a14_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a13_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a12_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a10_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a9_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a7_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a6_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a4_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a3_a_aq,
fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a1_a_aq,fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout,fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout,
fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.ax_width = 24;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.ay_scan_in_width = 26;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.operation_mode = "m27x27";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.result_a_width = 50;
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.signed_max = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_DSP0.use_chainadder = "false";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.first_bit_number = 23;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama23";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai401_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_lcell_comb fp_functions_0_aadd_15_a36(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a36_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_15_a36.extended_lut = "off";
defparam fp_functions_0_aadd_15_a36.lut_mask = 64'h0000000000005555;
defparam fp_functions_0_aadd_15_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_16_a166(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpR_uid48_fpDivTest_o_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_16_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_16_a166_sumout),
	.cout(fp_functions_0_aadd_16_a167),
	.shareout());
defparam fp_functions_0_aadd_16_a166.extended_lut = "off";
defparam fp_functions_0_aadd_16_a166.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_16_a166.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_17_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a166_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a17.extended_lut = "off";
defparam fp_functions_0_aadd_17_a17.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_17_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a166_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a17.extended_lut = "off";
defparam fp_functions_0_aadd_18_a17.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a17.shared_arith = "off";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_bit_number = 15;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama15";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_bit_number = 16;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama16";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_bit_number = 17;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama17";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_bit_number = 18;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama18";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_bit_number = 19;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama19";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_bit_number = 20;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama20";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_bit_number = 21;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama21";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.address_width = 3;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.data_width = 1;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_address = 0;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_bit_number = 22;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.init_file = "none";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.last_address = 4;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_depth = 5;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_name = "fp_functions_0|redist6_loadded_uid58_fpdivtest_q_6_mem_dmem|auto_generated|altera_syncram_impl1|lutrama22";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_width = 24;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai2307_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_8_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_15_a41(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_15_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_15_a41_sumout),
	.cout(fp_functions_0_aadd_15_a42),
	.shareout());
defparam fp_functions_0_aadd_15_a41.extended_lut = "off";
defparam fp_functions_0_aadd_15_a41.lut_mask = 64'h0000000000005555;
defparam fp_functions_0_aadd_15_a41.shared_arith = "off";

fourteennm_ff fp_functions_0_aexpR_uid48_fpDivTest_o_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_15_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpR_uid48_fpDivTest_o_a8_a_aq));
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpR_uid48_fpDivTest_o_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_17_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a151_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a22.extended_lut = "off";
defparam fp_functions_0_aadd_17_a22.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_17_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a151_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a22.extended_lut = "off";
defparam fp_functions_0_aadd_18_a22.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a22.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_20_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid25_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a23_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a24_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a25_a_aq));
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai413_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai413_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai413_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 5;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 20;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 21;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist12_expxmy_uid47_fpdivtest_q_23_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 9;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_lcell_comb fp_functions_0_aadd_17_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a146_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a27.extended_lut = "off";
defparam fp_functions_0_aadd_17_a27.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_17_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a146_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a27.extended_lut = "off";
defparam fp_functions_0_aadd_18_a27.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a27.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_13_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai2329_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai2329_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai2329_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a0_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracXIsZero_uid25_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_4_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid25_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid25_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid25_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_11_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a132_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a1_sumout),
	.cout(fp_functions_0_aadd_11_a2),
	.shareout());
defparam fp_functions_0_aadd_11_a1.extended_lut = "off";
defparam fp_functions_0_aadd_11_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a6_sumout),
	.cout(fp_functions_0_aadd_11_a7),
	.shareout());
defparam fp_functions_0_aadd_11_a6.extended_lut = "off";
defparam fp_functions_0_aadd_11_a6.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a11_sumout),
	.cout(fp_functions_0_aadd_11_a12),
	.shareout());
defparam fp_functions_0_aadd_11_a11.extended_lut = "off";
defparam fp_functions_0_aadd_11_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a16_sumout),
	.cout(fp_functions_0_aadd_11_a17),
	.shareout());
defparam fp_functions_0_aadd_11_a16.extended_lut = "off";
defparam fp_functions_0_aadd_11_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a21_sumout),
	.cout(fp_functions_0_aadd_11_a22),
	.shareout());
defparam fp_functions_0_aadd_11_a21.extended_lut = "off";
defparam fp_functions_0_aadd_11_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a26_sumout),
	.cout(fp_functions_0_aadd_11_a27),
	.shareout());
defparam fp_functions_0_aadd_11_a26.extended_lut = "off";
defparam fp_functions_0_aadd_11_a26.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a31_sumout),
	.cout(fp_functions_0_aadd_11_a32),
	.shareout());
defparam fp_functions_0_aadd_11_a31.extended_lut = "off";
defparam fp_functions_0_aadd_11_a31.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a36_sumout),
	.cout(fp_functions_0_aadd_11_a37),
	.shareout());
defparam fp_functions_0_aadd_11_a36.extended_lut = "off";
defparam fp_functions_0_aadd_11_a36.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a41_sumout),
	.cout(fp_functions_0_aadd_11_a42),
	.shareout());
defparam fp_functions_0_aadd_11_a41.extended_lut = "off";
defparam fp_functions_0_aadd_11_a41.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a46_sumout),
	.cout(fp_functions_0_aadd_11_a47),
	.shareout());
defparam fp_functions_0_aadd_11_a46.extended_lut = "off";
defparam fp_functions_0_aadd_11_a46.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a51_sumout),
	.cout(fp_functions_0_aadd_11_a52),
	.shareout());
defparam fp_functions_0_aadd_11_a51.extended_lut = "off";
defparam fp_functions_0_aadd_11_a51.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a56_sumout),
	.cout(fp_functions_0_aadd_11_a57),
	.shareout());
defparam fp_functions_0_aadd_11_a56.extended_lut = "off";
defparam fp_functions_0_aadd_11_a56.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a61_sumout),
	.cout(fp_functions_0_aadd_11_a62),
	.shareout());
defparam fp_functions_0_aadd_11_a61.extended_lut = "off";
defparam fp_functions_0_aadd_11_a61.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a66_sumout),
	.cout(fp_functions_0_aadd_11_a67),
	.shareout());
defparam fp_functions_0_aadd_11_a66.extended_lut = "off";
defparam fp_functions_0_aadd_11_a66.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a71_sumout),
	.cout(fp_functions_0_aadd_11_a72),
	.shareout());
defparam fp_functions_0_aadd_11_a71.extended_lut = "off";
defparam fp_functions_0_aadd_11_a71.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a76_sumout),
	.cout(fp_functions_0_aadd_11_a77),
	.shareout());
defparam fp_functions_0_aadd_11_a76.extended_lut = "off";
defparam fp_functions_0_aadd_11_a76.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a81_sumout),
	.cout(fp_functions_0_aadd_11_a82),
	.shareout());
defparam fp_functions_0_aadd_11_a81.extended_lut = "off";
defparam fp_functions_0_aadd_11_a81.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a86_sumout),
	.cout(fp_functions_0_aadd_11_a87),
	.shareout());
defparam fp_functions_0_aadd_11_a86.extended_lut = "off";
defparam fp_functions_0_aadd_11_a86.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a91_sumout),
	.cout(fp_functions_0_aadd_11_a92),
	.shareout());
defparam fp_functions_0_aadd_11_a91.extended_lut = "off";
defparam fp_functions_0_aadd_11_a91.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a96(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a96_sumout),
	.cout(fp_functions_0_aadd_11_a97),
	.shareout());
defparam fp_functions_0_aadd_11_a96.extended_lut = "off";
defparam fp_functions_0_aadd_11_a96.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a101(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a101_sumout),
	.cout(fp_functions_0_aadd_11_a102),
	.shareout());
defparam fp_functions_0_aadd_11_a101.extended_lut = "off";
defparam fp_functions_0_aadd_11_a101.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a106(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a106_sumout),
	.cout(fp_functions_0_aadd_11_a107),
	.shareout());
defparam fp_functions_0_aadd_11_a106.extended_lut = "off";
defparam fp_functions_0_aadd_11_a106.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a111(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a111_sumout),
	.cout(fp_functions_0_aadd_11_a112),
	.shareout());
defparam fp_functions_0_aadd_11_a111.extended_lut = "off";
defparam fp_functions_0_aadd_11_a111.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a116(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a116_sumout),
	.cout(fp_functions_0_aadd_11_a117),
	.shareout());
defparam fp_functions_0_aadd_11_a116.extended_lut = "off";
defparam fp_functions_0_aadd_11_a116.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a116.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a121(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a121_sumout),
	.cout(fp_functions_0_aadd_11_a122),
	.shareout());
defparam fp_functions_0_aadd_11_a121.extended_lut = "off";
defparam fp_functions_0_aadd_11_a121.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a121.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a126(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a126_sumout),
	.cout(fp_functions_0_aadd_11_a127),
	.shareout());
defparam fp_functions_0_aadd_11_a126.extended_lut = "off";
defparam fp_functions_0_aadd_11_a126.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a126.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_9_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_17_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a141_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a32.extended_lut = "off";
defparam fp_functions_0_aadd_17_a32.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_17_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a141_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a32.extended_lut = "off";
defparam fp_functions_0_aadd_18_a32.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a32.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_18_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_14_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[23]),
	.datad(!a[23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a1_sumout),
	.cout(fp_functions_0_aadd_14_a2),
	.shareout());
defparam fp_functions_0_aadd_14_a1.extended_lut = "off";
defparam fp_functions_0_aadd_14_a1.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a1.shared_arith = "off";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a1_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a2_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a3_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a4_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a5_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a6_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a7_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracYPostZ_uid56_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai119_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_bit_number = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama15";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_bit_number = 16;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama16";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_bit_number = 17;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama17";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_bit_number = 18;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama18";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_bit_number = 19;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama19";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_bit_number = 20;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama20";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_bit_number = 21;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama21";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.address_width = 4;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.data_width = 1;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_address = 0;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_bit_number = 22;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.init_file = "none";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.last_address = 14;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_depth = 15;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_name = "fp_functions_0|redist25_fracx_uid10_fpdivtest_b_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama22";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_width = 23;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.mixed_port_feed_through_mode = "dont care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "26961295370EF468740C1ECEE2DA0836A169A08AEDB99A2FD80B7BBFB893B955EA3E54D7D56DD48DB89083330C8C1019E77F7A98856FF060FF0CB910F64CE8C8";

fourteennm_lcell_comb fp_functions_0_aadd_11_a132(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a137_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_11_a132_cout),
	.shareout());
defparam fp_functions_0_aadd_11_a132.extended_lut = "off";
defparam fp_functions_0_aadd_11_a132.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a132.shared_arith = "off";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "16BF71007A796F7B43F8C5AC233A5A3F3BF257000C571D5DCCAF0484848A38C1696BB63F8D7B8C6B2C4CE1111DB562DD37F12C58438B2CC4E69A3B08E3D706A8";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "0C9C96C456D0934A900520AB63F2A0D039CF10046AE5F2B43802FD4E7D4B6F04CBF3BF5C96E2F1E132428A9A96040018E03A99C2E9466EEB2245AF7D4F5F1DC4";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "0222F920A8536D64B003428B7A6E88B038848331ADF9F44A63760379304EE5DF1056C9FB32903BE558C1EA36FE2E321A701A2F033CD24C0E60421BF87845C204";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "0194F5E8441492EC1666B2FAA1A38D8FC7A85E1DA26794E25D04AA7A1DFF850442CE508E4292281C710C848E5C518619633E308F216014A42D944AFA1D1FBECC";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "AAD8F34FD7C7A167AC3C4A17AE50174CCCA9AD90170E9CA33E5266D3F62EEBDF5AF2F9C8EC6632A98A2D46B2FB117B4D94B059C86181755194182860EB37181C";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "002C3C1654FE0C04A4DB1E9217123BB4B4EC21642FA0CCC90064B49C0D4E4F624D8A70D46C62F002CA7FB053E84E56C4A79E8F2B7866BD11794AB6913E9468BC";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "4447B776BADC476A8071DA0049D51B1FE008F835ACF9703E99E15E866542E94DDC9EECAE54F3D2221B0BD0B3586ACE3C6D21AF499096E17D67F558392236F27C";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "282867265E62826497DF670BD0920CA2E84AEF4E72EF77BBA5C2235C3EFA6052180F3813F5352AFADDC183EA0B405865850CA9446C9570BA0EEEE88336220356";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "1AB012463481AB9DD8358153CAEEAF94E5764F2814E58D393C814162BD789A4BCFAEBAF424B212473085A11283041BC1BEB820523805C8E49393941BF7A2CF54";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "066AA479F25533FC4AA600C96CFE65271CD48F1AA71CA9C76900D5819679AC469064C65811315DD40AFCC0A2532833D6686F8F1EBAF1D042F45EF7A6192A7B10";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "01E66D2AA499C3FC3992AA9270FE1C92A9670F066D56CE00E4AA99FF8D2D3041B548FE3559CF3567F9A900689CE55C32B01ACF34C659CA81A7CB0D3EA08DD338";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "001E1CE66DB4A956AD24CCE380FE038E64D2A5AB4998F0001C664B5529B1C0407325AB599E00F32D52CE0019B5499FF195530F0DAB61C6553839563E6ACFC9A0";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "0001FC1E1C7398CD9B6DA5A955AB552B4964C9CC71E0FFFFFC1E38CC9B6B55155A49339E1FFFF0E3365AAAAD2671E00F8CC95A56CC7E3E336AAD983E19A56DC0";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "000003FE03F0783C78E39C6733993366DB2DA4A52B55AAAAA954AD692DB26666638E3C1FE0000FE0F1C6666492D4AAAAD6926C670F8001F0E664B56B52C98E00";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "AAAAAAAB555AAD56AD4AD6B5A52DA5B4924936C9B266CCCCCE67318E31C3878783F03FE00000001FF03E1E1C71CC66664DB6DAD2A555555AB4B6D9B39CF1F000";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "66666666CCC99B3264D9B26C9364936DB6DB6DA496D25A5A5AD294A56B56AD52A9556AAAAAAAAAAAA554AB56A5694B4B69249364C999999CC738E1C3E0FE0000";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "1E1E1E1E3C3878F1E3C78E1C70E38F1C71C71C638E31C639C6318C6318CE633198CCE666666666666CCD99326CDB26D92492492DA4B4B4B5AD6A54A955AAAAAA";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_bit_number = 21;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_bit_number = 21;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mem_init0 = "01FE01FE03F807F01FC07E03F01F80FC0FC0FC1F81F03E07C1F07C1F07C1E0F0783C1E1E1E1E1E1E1C3C78F1E3C71E38E38E38E39C738C739CE63398CC666666";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_bit_number = 22;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_bit_number = 22;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mem_init0 = "0001FFFE0007FFF0003FFE000FFF8003FFC003FF800FFE003FF003FF003FE00FF803FE01FE01FE01FC03F80FE03F01F81F81F81F83F07C0F83E1F0783C1E1E1E";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_bit_number = 23;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_bit_number = 23;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mem_init0 = "00000001FFFFFFF0000001FFFFFF8000003FFFFF800001FFFFF00000FFFFE00007FFFE0001FFFE0003FFF8001FFF0007FF8007FF800FFC007FE00FF803FE01FE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_bit_number = 24;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_bit_number = 24;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mem_init0 = "000000000000000FFFFFFFFFFFFF8000000000007FFFFFFFFFF0000000001FFFFFFFFE00000001FFFFFFF8000000FFFFFF8000007FFFFC00001FFFF80001FFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_bit_number = 25;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_bit_number = 25;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mem_init0 = "00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFF80000000000007FFFFFFFFFFC0000000007FFFFFFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_bit_number = 26;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_bit_number = 26;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mem_init0 = "000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_bit_number = 27;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_bit_number = 27;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_bit_number = 28;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_bit_number = 28;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

fourteennm_ff fp_functions_0_aexpXmY_uid47_fpDivTest_o_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_14_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a8_a_aq));
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXmY_uid47_fpDivTest_o_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_17_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a136_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a37.extended_lut = "off";
defparam fp_functions_0_aadd_17_a37.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_17_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a136_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a37.extended_lut = "off";
defparam fp_functions_0_aadd_18_a37.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_14_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_14_a7.extended_lut = "off";
defparam fp_functions_0_aadd_14_a7.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_14_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[24]),
	.datad(!a[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a11_sumout),
	.cout(fp_functions_0_aadd_14_a12),
	.shareout());
defparam fp_functions_0_aadd_14_a11.extended_lut = "off";
defparam fp_functions_0_aadd_14_a11.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[25]),
	.datad(!a[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a16_sumout),
	.cout(fp_functions_0_aadd_14_a17),
	.shareout());
defparam fp_functions_0_aadd_14_a16.extended_lut = "off";
defparam fp_functions_0_aadd_14_a16.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[26]),
	.datad(!a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a21_sumout),
	.cout(fp_functions_0_aadd_14_a22),
	.shareout());
defparam fp_functions_0_aadd_14_a21.extended_lut = "off";
defparam fp_functions_0_aadd_14_a21.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[27]),
	.datad(!a[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a26_sumout),
	.cout(fp_functions_0_aadd_14_a27),
	.shareout());
defparam fp_functions_0_aadd_14_a26.extended_lut = "off";
defparam fp_functions_0_aadd_14_a26.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[28]),
	.datad(!a[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a31_sumout),
	.cout(fp_functions_0_aadd_14_a32),
	.shareout());
defparam fp_functions_0_aadd_14_a31.extended_lut = "off";
defparam fp_functions_0_aadd_14_a31.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[29]),
	.datad(!a[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a36_sumout),
	.cout(fp_functions_0_aadd_14_a37),
	.shareout());
defparam fp_functions_0_aadd_14_a36.extended_lut = "off";
defparam fp_functions_0_aadd_14_a36.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[30]),
	.datad(!a[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a41_sumout),
	.cout(fp_functions_0_aadd_14_a42),
	.shareout());
defparam fp_functions_0_aadd_14_a41.extended_lut = "off";
defparam fp_functions_0_aadd_14_a41.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_14_a41.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracYPostZ_uid56_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_afracYPostZ_uid56_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracYPostZ_uid56_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracYPostZ_uid56_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_19_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a22_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a21_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a20_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a19_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a18_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a17_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a16_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a15_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a14_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a13_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a12_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a11_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a10_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a8_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a7_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a5_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a4_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a2_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a1_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a13_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a12_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a10_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a9_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a7_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a6_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a4_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a3_a_aq,
fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a1_a_aq,fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout,fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout,
fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.ax_width = 23;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.ay_scan_in_width = 14;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.operation_mode = "m27x27";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.result_a_width = 37;
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.signed_max = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "D1A7B71FFB419AD34780F5BDF89065539B7BEA5CDD33EDEE44F68CD9C322E59A47583B479A569AA84537ED7F30C57E3B4AF7A59CFC0E91DE6B20C62872DF0075";

fourteennm_lcell_comb fp_functions_0_aadd_11_a137(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a147_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_11_a137_cout),
	.shareout());
defparam fp_functions_0_aadd_11_a137.extended_lut = "off";
defparam fp_functions_0_aadd_11_a137.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a137.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_14_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_14_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_14_a46_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_14_a46.extended_lut = "off";
defparam fp_functions_0_aadd_14_a46.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_14_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_17_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a131_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a42.extended_lut = "off";
defparam fp_functions_0_aadd_17_a42.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_17_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a131_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a42.extended_lut = "off";
defparam fp_functions_0_aadd_18_a42.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a42.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_11_a141(
	.dataa(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a29_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a141_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_11_a141.extended_lut = "off";
defparam fp_functions_0_aadd_11_a141.lut_mask = 64'h00000000000055AA;
defparam fp_functions_0_aadd_11_a141.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai134_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai138_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai138_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai138_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "6E00213CED44CAC6F411228681514A6D6A91CCAF691B25EA86C2706AC07F69C6C01C889AB54FF6704E0482940524F0255E4372D0C61E3590E6B007A5C27A13D0";

fourteennm_lcell_comb fp_functions_0_aadd_11_a147(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_11_a147_cout),
	.shareout());
defparam fp_functions_0_aadd_11_a147.extended_lut = "off";
defparam fp_functions_0_aadd_11_a147.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a147.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_17_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a126_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_17_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a47.extended_lut = "off";
defparam fp_functions_0_aadd_17_a47.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_17_a47.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a126_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_18_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a47.extended_lut = "off";
defparam fp_functions_0_aadd_18_a47.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_18_a47.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_first_bit_number = 29;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_first_bit_number = 29;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_3_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_lowRangeB_uid126_invPolyEval_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_lowRangeB_uid126_invPolyEval_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist2_lowRangeB_uid126_invPolyEval_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_lowRangeB_uid126_invPolyEval_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a0_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a1_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a2_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a3_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a4_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a5_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a6_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a7_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a8_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a9_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a10_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a11_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a12_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a13_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a14_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a15_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a16_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a17_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a18_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a19_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a20_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a21_a_aq));
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a8_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a9_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a10_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a11_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a12_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a13_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1513_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist11_yaddr_uid51_fpdivtest_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 9;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a8_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a4_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a3_a_aq,
fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a2_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC0_uid112_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC0_uid112_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 9;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 511;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 31;
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid112_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "2910A108D6843ED139497F1BAA7821D4C6F25BCAFE778362C9C4A5CA0C3F7575A6529A1DC2FFBE34211350D8F9B4A38835BA7C5305ADC9CC7B999768B4722528";

fourteennm_lcell_comb fp_functions_0_aadd_17_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a121_sumout),
	.datad(!fp_functions_0_aadd_16_a116_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_17_a52_cout),
	.shareout());
defparam fp_functions_0_aadd_17_a52.extended_lut = "off";
defparam fp_functions_0_aadd_17_a52.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_17_a52.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_18_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_16_a121_sumout),
	.datad(!fp_functions_0_aadd_16_a116_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_18_a52_cout),
	.shareout());
defparam fp_functions_0_aadd_18_a52.extended_lut = "off";
defparam fp_functions_0_aadd_18_a52.lut_mask = 64'h00000000F0000FF0;
defparam fp_functions_0_aadd_18_a52.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_6_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a1_sumout),
	.cout(fp_functions_0_aadd_6_a2),
	.shareout());
defparam fp_functions_0_aadd_6_a1.extended_lut = "off";
defparam fp_functions_0_aadd_6_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a6_sumout),
	.cout(fp_functions_0_aadd_6_a7),
	.shareout());
defparam fp_functions_0_aadd_6_a6.extended_lut = "off";
defparam fp_functions_0_aadd_6_a6.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a11_sumout),
	.cout(fp_functions_0_aadd_6_a12),
	.shareout());
defparam fp_functions_0_aadd_6_a11.extended_lut = "off";
defparam fp_functions_0_aadd_6_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a16_sumout),
	.cout(fp_functions_0_aadd_6_a17),
	.shareout());
defparam fp_functions_0_aadd_6_a16.extended_lut = "off";
defparam fp_functions_0_aadd_6_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a21_sumout),
	.cout(fp_functions_0_aadd_6_a22),
	.shareout());
defparam fp_functions_0_aadd_6_a21.extended_lut = "off";
defparam fp_functions_0_aadd_6_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a26_sumout),
	.cout(fp_functions_0_aadd_6_a27),
	.shareout());
defparam fp_functions_0_aadd_6_a26.extended_lut = "off";
defparam fp_functions_0_aadd_6_a26.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a31_sumout),
	.cout(fp_functions_0_aadd_6_a32),
	.shareout());
defparam fp_functions_0_aadd_6_a31.extended_lut = "off";
defparam fp_functions_0_aadd_6_a31.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a36_sumout),
	.cout(fp_functions_0_aadd_6_a37),
	.shareout());
defparam fp_functions_0_aadd_6_a36.extended_lut = "off";
defparam fp_functions_0_aadd_6_a36.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a41_sumout),
	.cout(fp_functions_0_aadd_6_a42),
	.shareout());
defparam fp_functions_0_aadd_6_a41.extended_lut = "off";
defparam fp_functions_0_aadd_6_a41.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a46_sumout),
	.cout(fp_functions_0_aadd_6_a47),
	.shareout());
defparam fp_functions_0_aadd_6_a46.extended_lut = "off";
defparam fp_functions_0_aadd_6_a46.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a51_sumout),
	.cout(fp_functions_0_aadd_6_a52),
	.shareout());
defparam fp_functions_0_aadd_6_a51.extended_lut = "off";
defparam fp_functions_0_aadd_6_a51.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a56_sumout),
	.cout(fp_functions_0_aadd_6_a57),
	.shareout());
defparam fp_functions_0_aadd_6_a56.extended_lut = "off";
defparam fp_functions_0_aadd_6_a56.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a61(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a61_sumout),
	.cout(fp_functions_0_aadd_6_a62),
	.shareout());
defparam fp_functions_0_aadd_6_a61.extended_lut = "off";
defparam fp_functions_0_aadd_6_a61.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a66(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a66_sumout),
	.cout(fp_functions_0_aadd_6_a67),
	.shareout());
defparam fp_functions_0_aadd_6_a66.extended_lut = "off";
defparam fp_functions_0_aadd_6_a66.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a71(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a71_sumout),
	.cout(fp_functions_0_aadd_6_a72),
	.shareout());
defparam fp_functions_0_aadd_6_a71.extended_lut = "off";
defparam fp_functions_0_aadd_6_a71.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a76(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a76_sumout),
	.cout(fp_functions_0_aadd_6_a77),
	.shareout());
defparam fp_functions_0_aadd_6_a76.extended_lut = "off";
defparam fp_functions_0_aadd_6_a76.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a81(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a81_sumout),
	.cout(fp_functions_0_aadd_6_a82),
	.shareout());
defparam fp_functions_0_aadd_6_a81.extended_lut = "off";
defparam fp_functions_0_aadd_6_a81.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a86(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a86_sumout),
	.cout(fp_functions_0_aadd_6_a87),
	.shareout());
defparam fp_functions_0_aadd_6_a86.extended_lut = "off";
defparam fp_functions_0_aadd_6_a86.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a91(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a91_sumout),
	.cout(fp_functions_0_aadd_6_a92),
	.shareout());
defparam fp_functions_0_aadd_6_a91.extended_lut = "off";
defparam fp_functions_0_aadd_6_a91.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a96(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a96_sumout),
	.cout(fp_functions_0_aadd_6_a97),
	.shareout());
defparam fp_functions_0_aadd_6_a96.extended_lut = "off";
defparam fp_functions_0_aadd_6_a96.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a101(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a101_sumout),
	.cout(fp_functions_0_aadd_6_a102),
	.shareout());
defparam fp_functions_0_aadd_6_a101.extended_lut = "off";
defparam fp_functions_0_aadd_6_a101.lut_mask = 64'h0000000011116666;
defparam fp_functions_0_aadd_6_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a106(
	.dataa(!fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(!fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a106_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_6_a106.extended_lut = "off";
defparam fp_functions_0_aadd_6_a106.lut_mask = 64'h0000000000006666;
defparam fp_functions_0_aadd_6_a106.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_14_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout,fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout,
fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.ax_width = 12;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.ay_scan_in_width = 12;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.operation_mode = "m18x18_full";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.result_a_width = 24;
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.signed_max = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "2E1DAB5CF8DD433CB78A33C2905FC81FF4ACEBF70A9AE12EBCB3189594F584596A9D2F4FF1952EECE484607ACF15A96FAC13EC8D2AD0902EEDC27FBEF1DC3EA8";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "4CF2A83262068783D44E881BCD67CDDE8DEC815F2B85FE5C9F249ED19E7D0979EB792CE8AC80F24090C85340FC09937B87DC5705217B7521B5671084F8B17C07";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "5E6316D0F6BFC122161C2241B5F2ECA8378135412BB1B360B195121D5E4A97B19874A2C829EB2A020C3A63FAFF25A0DD5F7CFAF61EFED47E3A1B8F16A8D3DF1A";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "6A057CB0AED3E8C9E215C997D253518DCCDE849191AE865DAE9D995A59376ED3CF1017ECBC83BEE7CE9FB0C9CCFBDCA7D85F8EE5EE8BC7EB3FFC2B1D25F3AE60";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "735300DA611AA7F2AE19581AB066C12409BF2C1B7D1F2E6BB5989D22DD050A18184E85FB1E77E3F0B53DD21A1E23C48EFC2E37DD2835AB2A5999ABD5AD81B96E";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "7C65AA49E01CCAA99E1E6D498F84949C0ED563E2548034D846CB9E5621ACF34812C0D3F280AFC9FA797EB344BF62B98A145F7A126DD17791BC3C105D40395C02";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "7F86336D4AB5A66781E07192D5524C7C0F19B556CC7FC76D52479F9B549C0392B63F1AA980CAA7FCAB00D93F2AE32B8CB395034FBBE4FA82817E82D8F429BEF6";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "7FF83C718CD934B52AAAD4B64CCE3C03F01E399B695552DB31C0601C66D6A9498E001CCD2A599FFF3255B7003349678F254CFC6A9806A9832B00D62153CC80AE";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "7FFFC07E0F1E38C6333366DB696B56AAAAB56B4924CCCE38F03FFFE078E7326D2B554A5B66387FFFC39925AA96D8E0703996AAD987F8CD296700E4AB300ED59E";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "D555552AA54A95AD69692DB6DB26CD99998CE738E3C3C1F80FFFFFFF80F83C71CC666C924B52AAAAA94B6C998E381FFFC1E7336D2AAA5B671F00F8CDA55A4C7E";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "999999B3366CD9364DB24924924B692D2D294A52B56A9552AAAAAAAAAA556AD4A52D25B6D93666666738E38781F8000001F83C71CCCC924A55AA55A49339C3FE";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "E1E1E1C3C78F1E3871C38E38E38C71CE31CE739CC673199CCCCCCCCCCC99B366C9B64924925B4B4B4A52B52AD552AAAAAB556AD4A5A5B6D93366339C70F83FFE";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "FE01FE03F80FE03F81FC0FC0FC0F81F03E0F83E0F87C1E1F0F0F0F0F0F1E3C78F1C78E38E39C738C739CC633199CCCCCCD99B366C936DB6DA5B4A5295AAD5554";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "FFFE0003FFF0003FFE000FFF000FFE003FF003FF007FE01FF00FF00FF01FC07F01F80FC0FC1F83F07C1F07C3E1E0F0F0F1E1C3870E38E38E39C739CE63319998";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "FFFFFFFC0000003FFFFFF000000FFFFFC00003FFFF80001FFFF0000FFFE0007FFE000FFF001FFC007FE007FC01FF00FF01FE03F80FC0FC0FC1F83E0F83C1E1E0";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "FFFFFFFFFFFFFFC000000000000FFFFFFFFFFC000000001FFFFFFFF00000007FFFFFF000001FFFFF800007FFFE0000FFFE0003FFF000FFF001FFC00FFC01FE00";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000001FFFFFFFFFFFFFFF8000000000001FFFFFFFFFF800000000FFFFFFFC000000FFFFFE00000FFFFE0000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000001FFFFFFFFFFFFFFFFFFF00000000000000FFFFFFFFFFF000000000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC1_uid115_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fp_functions_0|memoryC1_uid115_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 9;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 511;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 21;
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid115_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1191_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 3;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 4;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 5;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fp_functions_0|redist9_ype_uid52_fpdivtest_b_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 14;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1525_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1525_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1525_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_12_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_15_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a0_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a1_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a2_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a3_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a4_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a5_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a6_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a7_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a8_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a9_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a10_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a11_a_aq));
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1203_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1203_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1203_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a0_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a1_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a1_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai899_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist10_yaddr_uid51_fpdivtest_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 9;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "138758D0451960851267F354EF19F92149A79DD88BD6A27F1184EFBA9CD54B961F66F85CD2956FC2D59E18EC4AFB5F638230AFD7A5AFDF842B9702260D8699D4";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "3EE530C82D7D48B3691C488CA6C7CB908693707D7CC5EAADC3037B14A0C89109653D5A6291FDD1EC1CD84046308AB067D2C8704AA1C3E3754B1C02D97C314B17";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "01E0F3381D075C8F0703C7BC9E3C388FAF70F3C4FBCC671FC89E2772604448BB13ED36D64B4B0B5AB74A2AEEAAAF52B5662ABB53390CF97A8B1C3C871F912042";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "001FF007FD00BC80FF003F837E03F87F80F00FC3F83C1F03C781E0F1E3C3C7870F1CF1CE38C738C6733919DD9999366CD06196F694A5ABD55E49542A56DA4D9B";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "00000FFFFD00037FFF00007FFE0007FF800FFFC007FC00FFC07FE00FE03FC07F00FC0FC1F83F07C1F0F8F83C7878F1E3CE1871CE739C6733393B3266CDB6DB49";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "0000000002FFFFFFFF00000001FFFFFF8000003FFFFC00003FFFE0001FFFC000FFFC003FF800FFC00FF807FC07F80FE03E07F03E0F83E0F0F8F8F1E1C38E38C7";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "000000000000000000FFFFFFFFFFFFFF800000000003FFFFFFFFE00000003FFFFFFC000007FFFFC00007FFFC0007FFE001FFF001FF801FF007F80FE03F81F83F";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000003FFFFFFFFFFC000000003FFFFFFE000000FFFFF80000FFFF8001FFF8007FF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000003FFFFFFFFFFFFFFFE000000000007FFFFFFFF80000007FFFFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "00000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(areset),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,b[22],b[21],b[20],b[19],b[18],b[17],b[16],b[15],b[14]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Div_altera_fp_functions_191_j5x7yay_memoryC2_uid118_invTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC2_uid118_invTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 9;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 511;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 512;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid118_invTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a2_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a3_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a4_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a5_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a6_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a7_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a8_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a9_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a10_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a11_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a12_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a13_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_13_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a0_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a1_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_1_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_10_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a16_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a16_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a2_a(
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a2_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a3_a(
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a3_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a4_a(
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a4_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a5_a(
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a5_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a6_a(
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a6_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a7_a(
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a7_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a8_a(
	.clk(clk),
	.d(b[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a8_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a9_a(
	.clk(clk),
	.d(b[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a9_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a10_a(
	.clk(clk),
	.d(b[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a10_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a11_a(
	.clk(clk),
	.d(b[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a11_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a12_a(
	.clk(clk),
	.d(b[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a12_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a13_a(
	.clk(clk),
	.d(b[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a13_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a0_a(
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a0_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a1_a(
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a1_a_aq));
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_delay_0_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai911_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai911_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai911_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a17_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a17_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_11_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a18_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a18_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a19_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a19_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a20_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a20_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a21_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a21_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a23_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a22_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcZ_x_uid23_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq));
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcZ_y_uid37_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexpXIsMax_uid38_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq));
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid39_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq));
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexpXIsMax_uid24_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a22_a_a0_a_aq));
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a23_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_asignR_uid46_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a23_a_a0_a_aq));
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a23_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a23_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcZ_x_uid23_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_7_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexcZ_x_uid23_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcZ_x_uid23_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcZ_x_uid23_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcZ_y_uid37_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_6_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexcZ_y_uid37_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcZ_y_uid37_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcZ_y_uid37_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXIsMax_uid38_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_1_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXIsMax_uid38_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexpXIsMax_uid38_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXIsMax_uid38_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracXIsZero_uid39_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_16_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid39_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid39_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid39_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXIsMax_uid24_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_5_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXIsMax_uid24_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexpXIsMax_uid24_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXIsMax_uid24_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracYZero_uid15_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_asignR_uid46_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_asignR_uid46_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_asignR_uid46_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_asignR_uid46_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracYZero_uid15_fpDivTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_16_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_afracYZero_uid15_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracYZero_uid15_fpDivTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracYZero_uid15_fpDivTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1(
	.dataa(!fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist19_excI_x_uid27_fpDivTest_q_1_q_a0_a_aq),
	.datac(!fp_functions_0_aexpOvf_uid84_fpDivTest_o_a12_a_aq),
	.datad(!fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aredist17_excZ_y_uid37_fpDivTest_q_25_q_a0_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1.extended_lut = "off";
defparam fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1.lut_mask = 64'hEEAECC00EEAECC00;
defparam fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_31_a0(
	.dataa(!fp_functions_0_aexcR_y_uid45_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist18_excR_x_uid31_fpDivTest_q_1_q_a0_a_aq),
	.datac(!fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist23_excZ_x_uid23_fpDivTest_q_25_q_a0_a_aq),
	.datae(!fp_functions_0_aexpUdf_uid81_fpDivTest_o_a12_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_31_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_31_a0.extended_lut = "off";
defparam fp_functions_0_aMux_31_a0.lut_mask = 64'hE0A0F0A0E0A0F0A0;
defparam fp_functions_0_aMux_31_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_32_a2(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_32_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_32_a2.extended_lut = "off";
defparam fp_functions_0_aMux_32_a2.lut_mask = 64'h0007000700070007;
defparam fp_functions_0_aMux_32_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_31_a1(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_31_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_31_a1.extended_lut = "off";
defparam fp_functions_0_aMux_31_a1.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_31_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_30_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a2_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_30_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_30_a0.extended_lut = "off";
defparam fp_functions_0_aMux_30_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_30_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_29_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a3_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_29_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_29_a0.extended_lut = "off";
defparam fp_functions_0_aMux_29_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_29_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_28_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_28_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_28_a0.extended_lut = "off";
defparam fp_functions_0_aMux_28_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_28_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_27_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a5_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_27_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_27_a0.extended_lut = "off";
defparam fp_functions_0_aMux_27_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_27_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_26_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a6_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_26_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_26_a0.extended_lut = "off";
defparam fp_functions_0_aMux_26_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_26_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_25_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a7_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_25_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_25_a0.extended_lut = "off";
defparam fp_functions_0_aMux_25_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_25_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_24_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a8_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_24_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_24_a0.extended_lut = "off";
defparam fp_functions_0_aMux_24_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_24_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_23_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a9_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_23_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_23_a0.extended_lut = "off";
defparam fp_functions_0_aMux_23_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_23_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_22_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a10_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_22_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_22_a0.extended_lut = "off";
defparam fp_functions_0_aMux_22_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_22_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_21_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a11_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_21_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_21_a0.extended_lut = "off";
defparam fp_functions_0_aMux_21_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_21_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_20_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a12_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_20_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_20_a0.extended_lut = "off";
defparam fp_functions_0_aMux_20_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_20_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_19_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a13_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_19_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_19_a0.extended_lut = "off";
defparam fp_functions_0_aMux_19_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_19_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_18_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a14_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_18_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_18_a0.extended_lut = "off";
defparam fp_functions_0_aMux_18_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_18_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_17_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a15_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_17_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_17_a0.extended_lut = "off";
defparam fp_functions_0_aMux_17_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_17_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_16_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a16_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_16_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_16_a0.extended_lut = "off";
defparam fp_functions_0_aMux_16_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_16_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_15_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a17_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_15_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_15_a0.extended_lut = "off";
defparam fp_functions_0_aMux_15_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_15_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_14_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a18_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_14_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_14_a0.extended_lut = "off";
defparam fp_functions_0_aMux_14_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_14_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_13_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a19_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_13_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_13_a0.extended_lut = "off";
defparam fp_functions_0_aMux_13_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_13_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_12_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a20_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_12_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_12_a0.extended_lut = "off";
defparam fp_functions_0_aMux_12_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_12_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_11_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a21_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_11_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_11_a0.extended_lut = "off";
defparam fp_functions_0_aMux_11_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_11_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_10_a0(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist4_fracRPreExc_uid78_fpDivTest_b_1_q_a22_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_10_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_10_a0.extended_lut = "off";
defparam fp_functions_0_aMux_10_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_10_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a2(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a2.extended_lut = "off";
defparam fp_functions_0_aMux_9_a2.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a3(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a3.extended_lut = "off";
defparam fp_functions_0_aMux_9_a3.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a4(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a2_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a4.extended_lut = "off";
defparam fp_functions_0_aMux_9_a4.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a5(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a3_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a5.extended_lut = "off";
defparam fp_functions_0_aMux_9_a5.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a6(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a6.extended_lut = "off";
defparam fp_functions_0_aMux_9_a6.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a7(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a5_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a7.extended_lut = "off";
defparam fp_functions_0_aMux_9_a7.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a8(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a6_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a8.extended_lut = "off";
defparam fp_functions_0_aMux_9_a8.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a9(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist3_excRPreExc_uid79_fpDivTest_b_1_q_a7_a_aq),
	.datac(!fp_functions_0_aconcExc_uid98_fpDivTest_q_a1_a_a1_combout),
	.datad(!fp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a9.extended_lut = "off";
defparam fp_functions_0_aMux_9_a9.lut_mask = 64'h00A700A700A700A7;
defparam fp_functions_0_aMux_9_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_adivR_uid110_fpDivTest_q_a31_a(
	.dataa(!fp_functions_0_aexcRNaN_uid97_fpDivTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist13_signR_uid46_fpDivTest_q_25_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_adivR_uid110_fpDivTest_q_a31_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_adivR_uid110_fpDivTest_q_a31_a.extended_lut = "off";
defparam fp_functions_0_adivR_uid110_fpDivTest_q_a31_a.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_adivR_uid110_fpDivTest_q_a31_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1(
	.dataa(!fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datae(!fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1.lut_mask = 64'h1F11FFFF1F111F1F;
defparam fp_functions_0_aexcRNaN_uid97_fpDivTest_qi_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a9_a_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a(
	.dataa(!fp_functions_0_aredist16_excZ_y_uid37_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_aexcR_y_uid45_fpDivTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a(
	.dataa(!fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist20_fracXIsZero_uid25_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aexcI_x_uid27_fpDivTest_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a(
	.dataa(!fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_aexcR_x_uid31_fpDivTest_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0(
	.dataa(!fp_functions_0_aredist22_excZ_x_uid23_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist15_expXIsMax_uid38_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_aredist14_fracXIsZero_uid39_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist21_expXIsMax_uid24_fpDivTest_q_24_adelay_signals_a0_a_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0.lut_mask = 64'h0301030103010301;
defparam fp_functions_0_aregOrZeroOverInf_uid88_fpDivTest_qi_a0_a_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a49_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2642_a0(
	.dataa(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a_aq),
	.datad(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2642_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2642_a0.extended_lut = "off";
defparam fp_functions_0_ai2642_a0.lut_mask = 64'h02A202A202A202A2;
defparam fp_functions_0_ai2642_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2642_a1(
	.dataa(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq),
	.datae(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.dataf(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2642_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2642_a1.extended_lut = "off";
defparam fp_functions_0_ai2642_a1.lut_mask = 64'h20202A2A20752A7F;
defparam fp_functions_0_ai2642_a1.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0(
	.dataa(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a49_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2690_a0(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a0.extended_lut = "off";
defparam fp_functions_0_ai2690_a0.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a1(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a1.extended_lut = "off";
defparam fp_functions_0_ai2690_a1.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a1.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a2(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a2.extended_lut = "off";
defparam fp_functions_0_ai2690_a2.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a3(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a3.extended_lut = "off";
defparam fp_functions_0_ai2690_a3.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a3.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a4(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a4.extended_lut = "off";
defparam fp_functions_0_ai2690_a4.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a4.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a5(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a5.extended_lut = "off";
defparam fp_functions_0_ai2690_a5.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a5.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a6(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a6.extended_lut = "off";
defparam fp_functions_0_ai2690_a6.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a6.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a7(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a7.extended_lut = "off";
defparam fp_functions_0_ai2690_a7.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a7.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a8(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a8.extended_lut = "off";
defparam fp_functions_0_ai2690_a8.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a8.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a36_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a9(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a9.extended_lut = "off";
defparam fp_functions_0_ai2690_a9.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a9.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a37_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a10(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a10.extended_lut = "off";
defparam fp_functions_0_ai2690_a10.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a10.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a38_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a11(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a37_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a11.extended_lut = "off";
defparam fp_functions_0_ai2690_a11.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a11.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a39_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a12(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a12.extended_lut = "off";
defparam fp_functions_0_ai2690_a12.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a12.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a40_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a13(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a39_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a13.extended_lut = "off";
defparam fp_functions_0_ai2690_a13.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a13.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a41_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a14(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a40_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a14.extended_lut = "off";
defparam fp_functions_0_ai2690_a14.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a14.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a42_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a15(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a41_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a15.extended_lut = "off";
defparam fp_functions_0_ai2690_a15.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a15.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a43_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a16(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a42_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a16.extended_lut = "off";
defparam fp_functions_0_ai2690_a16.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a16.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a44_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a17(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a17.extended_lut = "off";
defparam fp_functions_0_ai2690_a17.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a17.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a45_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a18(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a44_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a18.extended_lut = "off";
defparam fp_functions_0_ai2690_a18.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a18.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a46_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a19(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a45_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a19.extended_lut = "off";
defparam fp_functions_0_ai2690_a19.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a19.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a47_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a20(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a46_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a20.extended_lut = "off";
defparam fp_functions_0_ai2690_a20.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a20.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a48_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_s0_a48_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a48_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a48_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a48_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2690_a21(
	.dataa(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a47_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq),
	.datac(!fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_delay_adelay_signals_a0_a_a48_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq),
	.datae(!fp_functions_0_aredist7_fracYPostZ_uid56_fpDivTest_q_7_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_anorm_uid67_fpDivTest_b_a0_a_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2690_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2690_a21.extended_lut = "off";
defparam fp_functions_0_ai2690_a21.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_ai2690_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a23_a(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ch_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a24_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a24_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a25_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_invY_uid54_fpDivTest_merged_bit_select_b_1_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a25_a_aq));
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid137_prodDivPreNormProd_uid60_fpDivTest_cma_ah_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai456_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai401_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai401_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai401_a0.extended_lut = "off";
defparam fp_functions_0_ai401_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai401_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq));
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai2418_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai2418_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2307_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2307_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2307_a0.extended_lut = "off";
defparam fp_functions_0_ai2307_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai2307_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai456_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai456_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai456_a0.extended_lut = "off";
defparam fp_functions_0_ai456_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai456_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_8(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_8_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_8.extended_lut = "off";
defparam fp_functions_0_areduce_nor_8.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_8.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai2329_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2418_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2418_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2418_a0.extended_lut = "off";
defparam fp_functions_0_ai2418_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai2418_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a3_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2418_a1(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2418_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2418_a1.extended_lut = "off";
defparam fp_functions_0_ai2418_a1.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai2418_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_wraddr_q_a4_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_20(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a0_combout),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a1_combout),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a3_combout),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a2_combout),
	.datae(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_cmp_b_a0_a_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_20_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_20.extended_lut = "off";
defparam fp_functions_0_areduce_nor_20.lut_mask = 64'h0000100000001000;
defparam fp_functions_0_areduce_nor_20.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai413_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai413_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai413_a0.extended_lut = "off";
defparam fp_functions_0_ai413_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai413_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai413_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai413_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai413_a1.extended_lut = "off";
defparam fp_functions_0_ai413_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai413_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai413_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai413_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai413_a2.extended_lut = "off";
defparam fp_functions_0_ai413_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai413_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aexpXmY_uid47_fpDivTest_o_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai2329_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2329_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2329_a0.extended_lut = "off";
defparam fp_functions_0_ai2329_a0.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2329_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0.lut_mask = 64'h7575757575757575;
defparam fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_13_a0(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_13_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_13_a0.extended_lut = "off";
defparam fp_functions_0_aadd_13_a0.lut_mask = 64'h6666666666666666;
defparam fp_functions_0_aadd_13_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2329_a1(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2329_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2329_a1.extended_lut = "off";
defparam fp_functions_0_ai2329_a1.lut_mask = 64'h1EF01EF01EF01EF0;
defparam fp_functions_0_ai2329_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2329_a2(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a_aq),
	.datae(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2329_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2329_a2.extended_lut = "off";
defparam fp_functions_0_ai2329_a2.lut_mask = 64'h01FEF00F01FEF00F;
defparam fp_functions_0_ai2329_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2329_a3(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a_aq),
	.datae(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a_aq),
	.dataf(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_eq_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2329_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2329_a3.extended_lut = "off";
defparam fp_functions_0_ai2329_a3.lut_mask = 64'h0001FFFE0FFFF000;
defparam fp_functions_0_ai2329_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4_a0(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a0_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a1_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a13_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a14_a_aq),
	.datae(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a18_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_4_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4_a1(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a5_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a6_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a7_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4_a1.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_4_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4_a2(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a2_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a11_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a20_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a21_a_aq),
	.datae(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a22_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4_a2.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_4_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a12_a_aq),
	.datab(!fp_functions_0_areduce_nor_4_a0_combout),
	.datac(!fp_functions_0_areduce_nor_4_a1_combout),
	.datad(!fp_functions_0_areduce_nor_4_a2_combout),
	.datae(!fp_functions_0_areduce_nor_4_a3_combout),
	.dataf(!fp_functions_0_areduce_nor_4_a4_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4.lut_mask = 64'h0000000000000002;
defparam fp_functions_0_areduce_nor_4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a36_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_areduce_nor_9(
	.dataa(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist6_lOAdded_uid58_fpDivTest_q_6_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_9_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_9.extended_lut = "off";
defparam fp_functions_0_areduce_nor_9.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_18(
	.dataa(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a3_a_aq),
	.datae(!fp_functions_0_aredist12_expXmY_uid47_fpDivTest_q_23_rdcnt_i_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_18_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_18.extended_lut = "off";
defparam fp_functions_0_areduce_nor_18.lut_mask = 64'h0000100000001000;
defparam fp_functions_0_areduce_nor_18.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai182_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai182_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai182_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai119_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai119_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai119_a0.extended_lut = "off";
defparam fp_functions_0_ai119_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai119_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(a[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(a[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(a[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a(
	.clk(clk),
	.d(a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a(
	.clk(clk),
	.d(a[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a(
	.clk(clk),
	.d(a[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a(
	.clk(clk),
	.d(a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a(
	.clk(clk),
	.d(a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a(
	.clk(clk),
	.d(a[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a(
	.clk(clk),
	.d(a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a(
	.clk(clk),
	.d(a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq));
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a(
	.dataa(!fp_functions_0_aredist24_fracYZero_uid15_fpDivTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aadd_11_a141_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_afracYPostZ_uid56_fpDivTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai182_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai182_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai182_a0.extended_lut = "off";
defparam fp_functions_0_ai182_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai182_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai182_a1(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai182_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai182_a1.extended_lut = "off";
defparam fp_functions_0_ai182_a1.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai182_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai182_a2(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai182_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai182_a2.extended_lut = "off";
defparam fp_functions_0_ai182_a2.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai182_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_wraddr_q_a3_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_19(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a0_combout),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a1_combout),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a2_combout),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_cmp_b_a0_a_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_19_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_19.extended_lut = "off";
defparam fp_functions_0_areduce_nor_19.lut_mask = 64'h0004000400040004;
defparam fp_functions_0_areduce_nor_19.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_lowRangeB_uid126_invPolyEval_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid128_invPolyEval_o_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ch_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai134_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai134_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai134_a0.extended_lut = "off";
defparam fp_functions_0_ai134_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai134_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai138_a0(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai138_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai138_a0.extended_lut = "off";
defparam fp_functions_0_ai138_a0.lut_mask = 64'h6C6C6C6C6C6C6C6C;
defparam fp_functions_0_ai138_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai138_a1(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai138_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai138_a1.extended_lut = "off";
defparam fp_functions_0_ai138_a1.lut_mask = 64'h1E3C1E3C1E3C1E3C;
defparam fp_functions_0_ai138_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai138_a2(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a_aq),
	.datae(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai138_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai138_a2.extended_lut = "off";
defparam fp_functions_0_ai138_a2.lut_mask = 64'h01FE03FC01FE03FC;
defparam fp_functions_0_ai138_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid143_pT2_uid131_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_areduce_nor_3(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_rdcnt_i_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_3_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_3.lut_mask = 64'h0004000400040004;
defparam fp_functions_0_areduce_nor_3.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1544_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1513_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1513_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1513_a0.extended_lut = "off";
defparam fp_functions_0_ai1513_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai1513_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1544_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1544_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1544_a0.extended_lut = "off";
defparam fp_functions_0_ai1544_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai1544_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_14(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_14_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_14.extended_lut = "off";
defparam fp_functions_0_areduce_nor_14.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_14.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_memoryC2_uid118_invTables_lutmem_r_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid140_pT1_uid125_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1222_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1191_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1191_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1191_a0.extended_lut = "off";
defparam fp_functions_0_ai1191_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai1191_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_yPE_uid52_fpDivTest_b_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1525_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1525_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1525_a0.extended_lut = "off";
defparam fp_functions_0_ai1525_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai1525_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1525_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1525_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1525_a1.extended_lut = "off";
defparam fp_functions_0_ai1525_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai1525_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1525_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1525_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1525_a2.extended_lut = "off";
defparam fp_functions_0_ai1525_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai1525_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1222_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1222_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1222_a0.extended_lut = "off";
defparam fp_functions_0_ai1222_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai1222_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_12(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_12_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_12.extended_lut = "off";
defparam fp_functions_0_areduce_nor_12.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_15(
	.dataa(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist11_yAddr_uid51_fpDivTest_b_14_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_15_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_15.extended_lut = "off";
defparam fp_functions_0_areduce_nor_15.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1203_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1203_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1203_a0.extended_lut = "off";
defparam fp_functions_0_ai1203_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai1203_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1203_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1203_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1203_a1.extended_lut = "off";
defparam fp_functions_0_ai1203_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai1203_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1203_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1203_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1203_a2.extended_lut = "off";
defparam fp_functions_0_ai1203_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai1203_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai930_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(b[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai899_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_sticky_ena_q_a0_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai899_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai899_a0.extended_lut = "off";
defparam fp_functions_0_ai899_a0.lut_mask = 64'h3737373737373737;
defparam fp_functions_0_ai899_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(b[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(b[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(b[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(b[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(b[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(b[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(b[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_areduce_nor_13(
	.dataa(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist9_yPE_uid52_fpDivTest_b_10_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_13_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_13.extended_lut = "off";
defparam fp_functions_0_areduce_nor_13.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a0_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a1_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai930_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq),
	.datad(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai930_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai930_a0.extended_lut = "off";
defparam fp_functions_0_ai930_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fp_functions_0_ai930_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_wraddr_q_a2_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a0_combout),
	.datae(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10.lut_mask = 64'h000000D8000000D8;
defparam fp_functions_0_areduce_nor_10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai911_a0(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai911_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai911_a0.extended_lut = "off";
defparam fp_functions_0_ai911_a0.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai911_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai911_a1(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai911_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai911_a1.extended_lut = "off";
defparam fp_functions_0_ai911_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fp_functions_0_ai911_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai911_a2(
	.dataa(!en[0]),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai911_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai911_a2.extended_lut = "off";
defparam fp_functions_0_ai911_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fp_functions_0_ai911_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11(
	.dataa(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist10_yAddr_uid51_fpDivTest_b_7_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_areduce_nor_11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_7_a0(
	.dataa(!a[23]),
	.datab(!a[24]),
	.datac(!a[25]),
	.datad(!a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_7_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_7_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_7_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_7_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_7(
	.dataa(!a[27]),
	.datab(!a[28]),
	.datac(!a[29]),
	.datad(!a[30]),
	.datae(!fp_functions_0_areduce_nor_7_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_7_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_7.extended_lut = "off";
defparam fp_functions_0_areduce_nor_7.lut_mask = 64'h0000800000008000;
defparam fp_functions_0_areduce_nor_7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6_a0(
	.dataa(!b[23]),
	.datab(!b[24]),
	.datac(!b[25]),
	.datad(!b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_6_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6(
	.dataa(!b[27]),
	.datab(!b[28]),
	.datac(!b[29]),
	.datad(!b[30]),
	.datae(!fp_functions_0_areduce_nor_6_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6.lut_mask = 64'h0000800000008000;
defparam fp_functions_0_areduce_nor_6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1_a0(
	.dataa(!b[23]),
	.datab(!b[24]),
	.datac(!b[25]),
	.datad(!b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1_a0.lut_mask = 64'h0001000100010001;
defparam fp_functions_0_areduce_nor_1_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1(
	.dataa(!b[27]),
	.datab(!b[28]),
	.datac(!b[29]),
	.datad(!b[30]),
	.datae(!fp_functions_0_areduce_nor_1_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1.lut_mask = 64'h0000000100000001;
defparam fp_functions_0_areduce_nor_1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_16_a0(
	.dataa(!b[2]),
	.datab(!b[3]),
	.datac(!b[4]),
	.datad(!b[0]),
	.datae(!b[1]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_16_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_16_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_16_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_16_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_16_a1(
	.dataa(!b[6]),
	.datab(!b[7]),
	.datac(!b[8]),
	.datad(!b[9]),
	.datae(!b[10]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_16_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_16_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_16_a1.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_16_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_16_a2(
	.dataa(!b[18]),
	.datab(!b[19]),
	.datac(!b[20]),
	.datad(!b[21]),
	.datae(!b[22]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_16_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_16_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_16_a2.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_16_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_16_a3(
	.dataa(!b[14]),
	.datab(!b[15]),
	.datac(!b[16]),
	.datad(!b[17]),
	.datae(!b[12]),
	.dataf(!b[13]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_16_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_16_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_16_a3.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_areduce_nor_16_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_16(
	.dataa(!b[5]),
	.datab(!b[11]),
	.datac(!fp_functions_0_areduce_nor_16_a0_combout),
	.datad(!fp_functions_0_areduce_nor_16_a1_combout),
	.datae(!fp_functions_0_areduce_nor_16_a2_combout),
	.dataf(!fp_functions_0_areduce_nor_16_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_16_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_16.extended_lut = "off";
defparam fp_functions_0_areduce_nor_16.lut_mask = 64'h0000000000000008;
defparam fp_functions_0_areduce_nor_16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_5_a0(
	.dataa(!a[23]),
	.datab(!a[24]),
	.datac(!a[25]),
	.datad(!a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_5_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_5_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_5_a0.lut_mask = 64'h0001000100010001;
defparam fp_functions_0_areduce_nor_5_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_5(
	.dataa(!a[27]),
	.datab(!a[28]),
	.datac(!a[29]),
	.datad(!a[30]),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_5_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_5.extended_lut = "off";
defparam fp_functions_0_areduce_nor_5.lut_mask = 64'h0000000100000001;
defparam fp_functions_0_areduce_nor_5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a(
	.dataa(!a[31]),
	.datab(!b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a.lut_mask = 64'h6666666666666666;
defparam fp_functions_0_asignR_uid46_fpDivTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4_a3(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a9_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a10_a_aq),
	.datac(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a4_a_aq),
	.datad(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a15_a_aq),
	.datae(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a16_a_aq),
	.dataf(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a17_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4_a3.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_areduce_nor_4_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4_a4(
	.dataa(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a19_a_aq),
	.datab(!fp_functions_0_aredist25_fracX_uid10_fpDivTest_b_17_outputreg0_q_a3_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4_a4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4_a4.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_areduce_nor_4_a4.shared_arith = "off";

assign q[22] = fp_functions_0_aMux_10_a0_combout;

assign q[21] = fp_functions_0_aMux_11_a0_combout;

assign q[20] = fp_functions_0_aMux_12_a0_combout;

assign q[19] = fp_functions_0_aMux_13_a0_combout;

assign q[18] = fp_functions_0_aMux_14_a0_combout;

assign q[17] = fp_functions_0_aMux_15_a0_combout;

assign q[16] = fp_functions_0_aMux_16_a0_combout;

assign q[15] = fp_functions_0_aMux_17_a0_combout;

assign q[14] = fp_functions_0_aMux_18_a0_combout;

assign q[13] = fp_functions_0_aMux_19_a0_combout;

assign q[12] = fp_functions_0_aMux_20_a0_combout;

assign q[11] = fp_functions_0_aMux_21_a0_combout;

assign q[10] = fp_functions_0_aMux_22_a0_combout;

assign q[9] = fp_functions_0_aMux_23_a0_combout;

assign q[8] = fp_functions_0_aMux_24_a0_combout;

assign q[7] = fp_functions_0_aMux_25_a0_combout;

assign q[6] = fp_functions_0_aMux_26_a0_combout;

assign q[5] = fp_functions_0_aMux_27_a0_combout;

assign q[4] = fp_functions_0_aMux_28_a0_combout;

assign q[3] = fp_functions_0_aMux_29_a0_combout;

assign q[2] = fp_functions_0_aMux_30_a0_combout;

assign q[1] = fp_functions_0_aMux_31_a1_combout;

assign q[0] = fp_functions_0_aMux_32_a2_combout;

assign q[23] = fp_functions_0_aMux_9_a2_combout;

assign q[24] = fp_functions_0_aMux_9_a3_combout;

assign q[25] = fp_functions_0_aMux_9_a4_combout;

assign q[26] = fp_functions_0_aMux_9_a5_combout;

assign q[27] = fp_functions_0_aMux_9_a6_combout;

assign q[28] = fp_functions_0_aMux_9_a7_combout;

assign q[29] = fp_functions_0_aMux_9_a8_combout;

assign q[30] = fp_functions_0_aMux_9_a9_combout;

assign q[31] = fp_functions_0_adivR_uid110_fpDivTest_q_a31_a_acombout;

endmodule
