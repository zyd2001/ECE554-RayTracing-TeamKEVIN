// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/23/2021 00:22:30"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Float_Inv (
	q,
	clk,
	areset,
	a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	clk;
input 	areset;
input 	[31:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq;
wire fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a0_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a1_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a2_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a3_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a4_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a5_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a7_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a8_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a9_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a10_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a11_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a12_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a13_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a14_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a15_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a16_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a17_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a18_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a19_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a20_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a21_a_aq;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a22_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a0_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a1_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a2_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a3_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a4_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a5_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a6_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a7_a_aq;
wire fp_functions_0_asignR_uid57_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aadd_2_a1_sumout;
wire fp_functions_0_aadd_11_a1_sumout;
wire fp_functions_0_aadd_11_a2;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aadd_11_a6_sumout;
wire fp_functions_0_aadd_11_a7;
wire fp_functions_0_aadd_11_a11_sumout;
wire fp_functions_0_aadd_11_a12;
wire fp_functions_0_aadd_11_a16_sumout;
wire fp_functions_0_aadd_11_a17;
wire fp_functions_0_aadd_11_a21_sumout;
wire fp_functions_0_aadd_11_a22;
wire fp_functions_0_aadd_11_a26_sumout;
wire fp_functions_0_aadd_11_a27;
wire fp_functions_0_aadd_11_a31_sumout;
wire fp_functions_0_aadd_11_a32;
wire fp_functions_0_aadd_11_a36_sumout;
wire fp_functions_0_aadd_11_a37;
wire fp_functions_0_aadd_11_a41_sumout;
wire fp_functions_0_aadd_11_a42;
wire fp_functions_0_aadd_11_a46_sumout;
wire fp_functions_0_aadd_11_a47;
wire fp_functions_0_aadd_11_a51_sumout;
wire fp_functions_0_aadd_11_a52;
wire fp_functions_0_aadd_11_a56_sumout;
wire fp_functions_0_aadd_11_a57;
wire fp_functions_0_aadd_11_a61_sumout;
wire fp_functions_0_aadd_11_a62;
wire fp_functions_0_aadd_11_a66_sumout;
wire fp_functions_0_aadd_11_a67;
wire fp_functions_0_aadd_11_a71_sumout;
wire fp_functions_0_aadd_11_a72;
wire fp_functions_0_aadd_11_a76_sumout;
wire fp_functions_0_aadd_11_a77;
wire fp_functions_0_aadd_11_a81_sumout;
wire fp_functions_0_aadd_11_a82;
wire fp_functions_0_aadd_11_a86_sumout;
wire fp_functions_0_aadd_11_a87;
wire fp_functions_0_aadd_11_a91_sumout;
wire fp_functions_0_aadd_11_a92;
wire fp_functions_0_aadd_11_a96_sumout;
wire fp_functions_0_aadd_11_a97;
wire fp_functions_0_aadd_11_a101_sumout;
wire fp_functions_0_aadd_11_a102;
wire fp_functions_0_aadd_11_a106_sumout;
wire fp_functions_0_aadd_11_a107;
wire fp_functions_0_aadd_11_a111_sumout;
wire fp_functions_0_aadd_3_a1_sumout;
wire fp_functions_0_aadd_3_a2;
wire fp_functions_0_aadd_3_a6_sumout;
wire fp_functions_0_aadd_3_a7;
wire fp_functions_0_aadd_3_a11_sumout;
wire fp_functions_0_aadd_3_a12;
wire fp_functions_0_aadd_3_a16_sumout;
wire fp_functions_0_aadd_3_a17;
wire fp_functions_0_aadd_3_a21_sumout;
wire fp_functions_0_aadd_3_a22;
wire fp_functions_0_aadd_3_a26_sumout;
wire fp_functions_0_aadd_3_a27;
wire fp_functions_0_aadd_3_a31_sumout;
wire fp_functions_0_aadd_3_a32;
wire fp_functions_0_aadd_3_a36_sumout;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aadd_2_a6_sumout;
wire fp_functions_0_aadd_2_a7;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_aadd_11_a117_cout;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a;
wire fp_functions_0_aadd_3_a42_cout;
wire fp_functions_0_aadd_2_a11_sumout;
wire fp_functions_0_aadd_2_a12;
wire fp_functions_0_aadd_2_a16_sumout;
wire fp_functions_0_aadd_2_a17;
wire fp_functions_0_aadd_2_a21_sumout;
wire fp_functions_0_aadd_2_a22;
wire fp_functions_0_aadd_2_a26_sumout;
wire fp_functions_0_aadd_2_a27;
wire fp_functions_0_aadd_2_a31_sumout;
wire fp_functions_0_aadd_2_a32;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a24_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a25_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a26_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a27_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a28_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a29_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a30_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a31_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a32_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a33_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a34_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a35_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a36_a;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_aadd_11_a122_cout;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aadd_2_a37_cout;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_aadd_11_a127_cout;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aadd_2_a42_cout;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist5_lowRangeB_uid74_invPolyEval_b_1_q_a0_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a0_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a1_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a2_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a3_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a4_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a5_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a6_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a7_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a8_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a9_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a10_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a11_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a12_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a13_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a14_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a15_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a16_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a17_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a18_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a19_a_aq;
wire fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a20_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a8_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a9_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a10_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a11_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a12_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a13_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a14_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aadd_2_a47_cout;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aadd_6_a1_sumout;
wire fp_functions_0_aadd_6_a2;
wire fp_functions_0_aadd_6_a6_sumout;
wire fp_functions_0_aadd_6_a7;
wire fp_functions_0_aadd_6_a11_sumout;
wire fp_functions_0_aadd_6_a12;
wire fp_functions_0_aadd_6_a16_sumout;
wire fp_functions_0_aadd_6_a17;
wire fp_functions_0_aadd_6_a21_sumout;
wire fp_functions_0_aadd_6_a22;
wire fp_functions_0_aadd_6_a26_sumout;
wire fp_functions_0_aadd_6_a27;
wire fp_functions_0_aadd_6_a31_sumout;
wire fp_functions_0_aadd_6_a32;
wire fp_functions_0_aadd_6_a36_sumout;
wire fp_functions_0_aadd_6_a37;
wire fp_functions_0_aadd_6_a41_sumout;
wire fp_functions_0_aadd_6_a42;
wire fp_functions_0_aadd_6_a46_sumout;
wire fp_functions_0_aadd_6_a47;
wire fp_functions_0_aadd_6_a51_sumout;
wire fp_functions_0_aadd_6_a52;
wire fp_functions_0_aadd_6_a56_sumout;
wire fp_functions_0_aadd_6_a57;
wire fp_functions_0_aadd_6_a61_sumout;
wire fp_functions_0_aadd_6_a62;
wire fp_functions_0_aadd_6_a66_sumout;
wire fp_functions_0_aadd_6_a67;
wire fp_functions_0_aadd_6_a71_sumout;
wire fp_functions_0_aadd_6_a72;
wire fp_functions_0_aadd_6_a76_sumout;
wire fp_functions_0_aadd_6_a77;
wire fp_functions_0_aadd_6_a81_sumout;
wire fp_functions_0_aadd_6_a82;
wire fp_functions_0_aadd_6_a86_sumout;
wire fp_functions_0_aadd_6_a87;
wire fp_functions_0_aadd_6_a91_sumout;
wire fp_functions_0_aadd_6_a92;
wire fp_functions_0_aadd_6_a96_sumout;
wire fp_functions_0_aadd_6_a97;
wire fp_functions_0_aadd_6_a101_sumout;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a0_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a1_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a2_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a3_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a4_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a5_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a6_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a7_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a8_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a9_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a10_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a11_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a12_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a13_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a14_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a15_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a16_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a17_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a18_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a19_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a20_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a21_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a22_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a23_a;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA24;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA25;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA26;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA27;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA28;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA29;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA30;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA31;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA32;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA33;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA34;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA35;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA36;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a7_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a0_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a1_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a2_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a3_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a4_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a5_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a6_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a7_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a8_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a9_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a10_a_aq;
wire fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a11_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a0_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a1_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a8_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a3_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a4_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a5_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a6_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a7_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a8_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a9_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a10_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a11_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a12_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a13_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a14_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a0_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a1_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a9_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a3_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a4_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a5_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a6_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a7_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a8_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a9_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a10_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a11_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a12_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a13_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a14_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a0_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a1_a_aq;
wire fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a10_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a11_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a12_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a13_a_a0_a_aq;
wire fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a14_a_a0_a_aq;
wire fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a15_a_a0_a_aq;
wire fp_functions_0_aMux_32_a2_combout;
wire fp_functions_0_aMux_31_a0_combout;
wire fp_functions_0_aMux_30_a0_combout;
wire fp_functions_0_aMux_29_a0_combout;
wire fp_functions_0_aMux_28_a0_combout;
wire fp_functions_0_aMux_27_a0_combout;
wire fp_functions_0_aMux_26_a0_combout;
wire fp_functions_0_aMux_25_a0_combout;
wire fp_functions_0_aMux_24_a0_combout;
wire fp_functions_0_aMux_23_a0_combout;
wire fp_functions_0_aMux_22_a0_combout;
wire fp_functions_0_aMux_21_a0_combout;
wire fp_functions_0_aMux_20_a0_combout;
wire fp_functions_0_aMux_19_a0_combout;
wire fp_functions_0_aMux_18_a0_combout;
wire fp_functions_0_aMux_17_a0_combout;
wire fp_functions_0_aMux_16_a0_combout;
wire fp_functions_0_aMux_15_a0_combout;
wire fp_functions_0_aMux_14_a0_combout;
wire fp_functions_0_aMux_13_a0_combout;
wire fp_functions_0_aMux_12_a0_combout;
wire fp_functions_0_aMux_11_a0_combout;
wire fp_functions_0_aMux_10_a0_combout;
wire fp_functions_0_aMux_9_a2_combout;
wire fp_functions_0_aMux_9_a3_combout;
wire fp_functions_0_aMux_9_a4_combout;
wire fp_functions_0_aMux_9_a5_combout;
wire fp_functions_0_aMux_9_a6_combout;
wire fp_functions_0_aMux_9_a7_combout;
wire fp_functions_0_aMux_9_a8_combout;
wire fp_functions_0_aMux_9_a9_combout;
wire fp_functions_0_areduce_nor_3_a0_combout;
wire fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a_acombout;
wire fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a_acombout;
wire fp_functions_0_areduce_nor_5_a0_combout;
wire fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0_combout;
wire fp_functions_0_areduce_nor_5_acombout;
wire fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout;
wire fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a_acombout;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq;
wire fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0_combout;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_cmpReg_q_a0_a_aq;
wire fp_functions_0_ai102_a0_combout;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fp_functions_0_ai138_a0_combout;
wire fp_functions_0_ai138_a1_combout;
wire fp_functions_0_ai138_a2_combout;
wire fp_functions_0_ai100_a0_combout;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq_aq;
wire fp_functions_0_ai112_a0_combout;
wire fp_functions_0_ai116_a0_combout;
wire fp_functions_0_ai116_a1_combout;
wire fp_functions_0_ai116_a2_combout;
wire fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_cmpReg_q_a0_a_aq;
wire fp_functions_0_ai1326_a0_combout;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fp_functions_0_ai1348_a0_combout;
wire fp_functions_0_ai1324_a0_combout;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_cmpReg_q_a0_a_aq;
wire fp_functions_0_ai1063_a0_combout;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq_aq;
wire fp_functions_0_ai1334_a0_combout;
wire fp_functions_0_ai1334_a1_combout;
wire fp_functions_0_ai1334_a2_combout;
wire fp_functions_0_ai1085_a0_combout;
wire fp_functions_0_ai1061_a0_combout;
wire fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq_aq;
wire fp_functions_0_ai1071_a0_combout;
wire fp_functions_0_ai1071_a1_combout;
wire fp_functions_0_ai1071_a2_combout;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_cmpReg_q_a0_a_aq;
wire fp_functions_0_ai825_a0_combout;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fp_functions_0_ai847_a0_combout;
wire fp_functions_0_ai823_a0_combout;
wire fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq_aq;
wire fp_functions_0_ai833_a0_combout;
wire fp_functions_0_ai833_a1_combout;
wire fp_functions_0_ai833_a2_combout;
wire fp_functions_0_afracXIsZero_uid23_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0_combout;
wire fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1_combout;
wire fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2_combout;
wire fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3_combout;
wire fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4_combout;

wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus;
wire [63:0] fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [63:0] fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus[0];

assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a0_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a1_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a2_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a3_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a4_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a5_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a6_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a7_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a8_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a9_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a10_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a11_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a12_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a13_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a14_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a15_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a16_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a17_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a18_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a19_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a20_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a21_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a22_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a23_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a24_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a25_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a26_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a27_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a28_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a29_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a30_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a31_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a32_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a33_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a34_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a35_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a36_a = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA37 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA38 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA39 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA40 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA41 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA42 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA43 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA44 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA45 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA46 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA47 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA48 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA49 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a0_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a1_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a2_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a3_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a4_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a5_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a6_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a7_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a8_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a9_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a10_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a11_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a12_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a13_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a14_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a15_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a16_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a17_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a18_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a19_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a20_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a21_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a22_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a23_a = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA24 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA25 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA26 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA27 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA28 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA29 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA30 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA31 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA32 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA33 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA34 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA35 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA36 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA37 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA38 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA39 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA40 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA41 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA42 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA43 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA44 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA45 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA46 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA47 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA48 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA49 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA50 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA51 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA52 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA53 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA54 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA55 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA56 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA57 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA58 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA59 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA60 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA61 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA62 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_aDATAOUTA63 = fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

fourteennm_ff fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_5_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a0_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a1_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a2_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a3_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a4_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a5_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a7_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a8_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a9_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a10_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a11_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a12_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a13_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a14_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a15_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a16_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a17_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a18_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a19_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a20_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a21_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_11_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a22_a_aq));
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a0_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a1_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a2_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a3_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a4_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a5_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a6_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a7_a_aq));
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_asignR_uid57_fpInverseTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_asignR_uid57_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_asignR_uid57_fpInverseTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_asignR_uid57_fpInverseTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a1.extended_lut = "off";
defparam fp_functions_0_aadd_2_a1.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_2_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a117_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a1_sumout),
	.cout(fp_functions_0_aadd_11_a2),
	.shareout());
defparam fp_functions_0_aadd_11_a1.extended_lut = "off";
defparam fp_functions_0_aadd_11_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a1.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_11_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a6_sumout),
	.cout(fp_functions_0_aadd_11_a7),
	.shareout());
defparam fp_functions_0_aadd_11_a6.extended_lut = "off";
defparam fp_functions_0_aadd_11_a6.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a11_sumout),
	.cout(fp_functions_0_aadd_11_a12),
	.shareout());
defparam fp_functions_0_aadd_11_a11.extended_lut = "off";
defparam fp_functions_0_aadd_11_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a16_sumout),
	.cout(fp_functions_0_aadd_11_a17),
	.shareout());
defparam fp_functions_0_aadd_11_a16.extended_lut = "off";
defparam fp_functions_0_aadd_11_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a21_sumout),
	.cout(fp_functions_0_aadd_11_a22),
	.shareout());
defparam fp_functions_0_aadd_11_a21.extended_lut = "off";
defparam fp_functions_0_aadd_11_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a26_sumout),
	.cout(fp_functions_0_aadd_11_a27),
	.shareout());
defparam fp_functions_0_aadd_11_a26.extended_lut = "off";
defparam fp_functions_0_aadd_11_a26.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a31_sumout),
	.cout(fp_functions_0_aadd_11_a32),
	.shareout());
defparam fp_functions_0_aadd_11_a31.extended_lut = "off";
defparam fp_functions_0_aadd_11_a31.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a36_sumout),
	.cout(fp_functions_0_aadd_11_a37),
	.shareout());
defparam fp_functions_0_aadd_11_a36.extended_lut = "off";
defparam fp_functions_0_aadd_11_a36.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a41_sumout),
	.cout(fp_functions_0_aadd_11_a42),
	.shareout());
defparam fp_functions_0_aadd_11_a41.extended_lut = "off";
defparam fp_functions_0_aadd_11_a41.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a46_sumout),
	.cout(fp_functions_0_aadd_11_a47),
	.shareout());
defparam fp_functions_0_aadd_11_a46.extended_lut = "off";
defparam fp_functions_0_aadd_11_a46.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a51_sumout),
	.cout(fp_functions_0_aadd_11_a52),
	.shareout());
defparam fp_functions_0_aadd_11_a51.extended_lut = "off";
defparam fp_functions_0_aadd_11_a51.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a56_sumout),
	.cout(fp_functions_0_aadd_11_a57),
	.shareout());
defparam fp_functions_0_aadd_11_a56.extended_lut = "off";
defparam fp_functions_0_aadd_11_a56.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a61_sumout),
	.cout(fp_functions_0_aadd_11_a62),
	.shareout());
defparam fp_functions_0_aadd_11_a61.extended_lut = "off";
defparam fp_functions_0_aadd_11_a61.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a66_sumout),
	.cout(fp_functions_0_aadd_11_a67),
	.shareout());
defparam fp_functions_0_aadd_11_a66.extended_lut = "off";
defparam fp_functions_0_aadd_11_a66.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a71_sumout),
	.cout(fp_functions_0_aadd_11_a72),
	.shareout());
defparam fp_functions_0_aadd_11_a71.extended_lut = "off";
defparam fp_functions_0_aadd_11_a71.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a76_sumout),
	.cout(fp_functions_0_aadd_11_a77),
	.shareout());
defparam fp_functions_0_aadd_11_a76.extended_lut = "off";
defparam fp_functions_0_aadd_11_a76.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a81_sumout),
	.cout(fp_functions_0_aadd_11_a82),
	.shareout());
defparam fp_functions_0_aadd_11_a81.extended_lut = "off";
defparam fp_functions_0_aadd_11_a81.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a86(
	.dataa(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a86_sumout),
	.cout(fp_functions_0_aadd_11_a87),
	.shareout());
defparam fp_functions_0_aadd_11_a86.extended_lut = "off";
defparam fp_functions_0_aadd_11_a86.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a91(
	.dataa(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a91_sumout),
	.cout(fp_functions_0_aadd_11_a92),
	.shareout());
defparam fp_functions_0_aadd_11_a91.extended_lut = "off";
defparam fp_functions_0_aadd_11_a91.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a96(
	.dataa(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a96_sumout),
	.cout(fp_functions_0_aadd_11_a97),
	.shareout());
defparam fp_functions_0_aadd_11_a96.extended_lut = "off";
defparam fp_functions_0_aadd_11_a96.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a101(
	.dataa(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a101_sumout),
	.cout(fp_functions_0_aadd_11_a102),
	.shareout());
defparam fp_functions_0_aadd_11_a101.extended_lut = "off";
defparam fp_functions_0_aadd_11_a101.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a106(
	.dataa(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a106_sumout),
	.cout(fp_functions_0_aadd_11_a107),
	.shareout());
defparam fp_functions_0_aadd_11_a106.extended_lut = "off";
defparam fp_functions_0_aadd_11_a106.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_11_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_11_a111(
	.dataa(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_11_a111_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_11_a111.extended_lut = "off";
defparam fp_functions_0_aadd_11_a111.lut_mask = 64'h00000000000055AA;
defparam fp_functions_0_aadd_11_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a1(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.datab(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a1_sumout),
	.cout(fp_functions_0_aadd_3_a2),
	.shareout());
defparam fp_functions_0_aadd_3_a1.extended_lut = "off";
defparam fp_functions_0_aadd_3_a1.lut_mask = 64'h0000000088886666;
defparam fp_functions_0_aadd_3_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a6(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0_combout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a6_sumout),
	.cout(fp_functions_0_aadd_3_a7),
	.shareout());
defparam fp_functions_0_aadd_3_a6.extended_lut = "off";
defparam fp_functions_0_aadd_3_a6.lut_mask = 64'h000000000F0AF0A5;
defparam fp_functions_0_aadd_3_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a11(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_2_a11_sumout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a11_sumout),
	.cout(fp_functions_0_aadd_3_a12),
	.shareout());
defparam fp_functions_0_aadd_3_a11.extended_lut = "off";
defparam fp_functions_0_aadd_3_a11.lut_mask = 64'h000000005F0AA0F5;
defparam fp_functions_0_aadd_3_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a16(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_2_a16_sumout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a16_sumout),
	.cout(fp_functions_0_aadd_3_a17),
	.shareout());
defparam fp_functions_0_aadd_3_a16.extended_lut = "off";
defparam fp_functions_0_aadd_3_a16.lut_mask = 64'h000000005F0AA0F5;
defparam fp_functions_0_aadd_3_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a21(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_2_a21_sumout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a21_sumout),
	.cout(fp_functions_0_aadd_3_a22),
	.shareout());
defparam fp_functions_0_aadd_3_a21.extended_lut = "off";
defparam fp_functions_0_aadd_3_a21.lut_mask = 64'h000000005F0AA0F5;
defparam fp_functions_0_aadd_3_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a26(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_2_a26_sumout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a26_sumout),
	.cout(fp_functions_0_aadd_3_a27),
	.shareout());
defparam fp_functions_0_aadd_3_a26.extended_lut = "off";
defparam fp_functions_0_aadd_3_a26.lut_mask = 64'h000000005F0AA0F5;
defparam fp_functions_0_aadd_3_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a31(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_2_a31_sumout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a31_sumout),
	.cout(fp_functions_0_aadd_3_a32),
	.shareout());
defparam fp_functions_0_aadd_3_a31.extended_lut = "off";
defparam fp_functions_0_aadd_3_a31.lut_mask = 64'h000000005F0AA0F5;
defparam fp_functions_0_aadd_3_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a36(
	.dataa(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_2_a6_sumout),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a36_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_3_a36.extended_lut = "off";
defparam fp_functions_0_aadd_3_a36.lut_mask = 64'h000000000000A0F5;
defparam fp_functions_0_aadd_3_a36.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai102_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 14;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 15;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist11_expx_uid6_fpinversetest_b_16_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a6_sumout),
	.cout(fp_functions_0_aadd_2_a7),
	.shareout());
defparam fp_functions_0_aadd_2_a6.extended_lut = "off";
defparam fp_functions_0_aadd_2_a6.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a6.shared_arith = "off";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "413A25F5D3B3988B07E2AEBDE3D8F9FB051955F86A911181F9740BA3AF6F307A";

fourteennm_lcell_comb fp_functions_0_aadd_11_a117(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a122_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_11_a117_cout),
	.shareout());
defparam fp_functions_0_aadd_11_a117.extended_lut = "off";
defparam fp_functions_0_aadd_11_a117.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a117.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "2690C5B24181CE001A153CAA9E3F4ABFD6FB6C5AC9828040C039FCAA884C4482";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "16B8AE426A4C1137F0E70A28F20C7F3282C68407D2268F2192431862369CFC6A";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "0C9BFB1326872C7AA13473216CADE29FC4D8AA4103A4B5DF60D891FD64089446";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "0226EE2A2D6474566A1A30E90A663AB8B8CEA8C08F4DCAEA3231CA75D8656586";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "AB3E4EB80DC09F5780C72DC659E2B89BE6A2EDC051C5C8A6B539469FBFC504CE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "00F2E80A7FB1C42088BACBF5381E6C8C4345F70CF91818CB321AA7C42A81621E";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "444A6117C71D8A36BEB06B3561987C49B24E244B43141259640C438A5565F0BE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "282DCF5E8209AEB36E34361B90F16D2A4AAC55FE0E80D05E8B364DC8EEF250D4";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "1AB0259E5404CE641B32BEA0A05F334978E7DB7BD1086BE444B6AD81393603D4";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "066AB61E32A90E12AC3194C06A9F1588D31D60D3CA05797D7D3319AF45E68B90";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "01E66D4B5B31F1F19A9AD8FFE64A59F7C9567FC96C032D8329CEAE65834653B8";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "001E1CC6C96B555AD3231F001E3934AA92678038DAAA4E00E4AB301CAA79C920";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "0001FC3E38E7333649694AAAAB5259331C780007C666DAAAB6CC3FFC66D56DC0";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "AAAAA954AD4A5A5B6DB26CCCCC639E3C1F8000003E1E3999925A9556B4998E00";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "666664CD9B26C936DB6925A5A5294A954AAAAAAAAB54AD2D2493266738E1F000";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "1E1E1C3C78E1C70E38E71C639CE7398CC666666666CD9B6492496D2D6A54AAAA";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "01FE03FC07E03F01F81F03E07C1F0783C1E1E1E1E1C3871C71C71CE319CC6666";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_bit_number = 21;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_bit_number = 21;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mem_init0 = "0001FFFC001FFF0007FF001FFC00FF803FE01FE01FC07F03F03F03E0F83C1E1E";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_bit_number = 22;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_bit_number = 22;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mem_init0 = "00000003FFFFFF000000FFFFFC00007FFFE0001FFFC000FFF000FFE007FC01FE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_bit_number = 23;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_bit_number = 23;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mem_init0 = "00000000000000FFFFFFFFFFFC000000001FFFFFFFC000000FFFFFE00003FFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_bit_number = 24;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_bit_number = 24;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mem_init0 = "00000000000000000000000003FFFFFFFFFFFFFFFFC000000000001FFFFFFFFE";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_bit_number = 25;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_bit_number = 25;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mem_init0 = "0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFE";

fourteennm_lcell_comb fp_functions_0_aadd_3_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a42.extended_lut = "off";
defparam fp_functions_0_aadd_3_a42.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_3_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a11_sumout),
	.cout(fp_functions_0_aadd_2_a12),
	.shareout());
defparam fp_functions_0_aadd_2_a11.extended_lut = "off";
defparam fp_functions_0_aadd_2_a11.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a16_sumout),
	.cout(fp_functions_0_aadd_2_a17),
	.shareout());
defparam fp_functions_0_aadd_2_a16.extended_lut = "off";
defparam fp_functions_0_aadd_2_a16.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a21_sumout),
	.cout(fp_functions_0_aadd_2_a22),
	.shareout());
defparam fp_functions_0_aadd_2_a21.extended_lut = "off";
defparam fp_functions_0_aadd_2_a21.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a26_sumout),
	.cout(fp_functions_0_aadd_2_a27),
	.shareout());
defparam fp_functions_0_aadd_2_a26.extended_lut = "off";
defparam fp_functions_0_aadd_2_a26.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a31_sumout),
	.cout(fp_functions_0_aadd_2_a32),
	.shareout());
defparam fp_functions_0_aadd_2_a31.extended_lut = "off";
defparam fp_functions_0_aadd_2_a31.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a31.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a21_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a20_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a19_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a18_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a17_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a16_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a15_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a14_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a13_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a12_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a14_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a13_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a12_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a10_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a9_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a7_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a6_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a4_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a3_a_aq,
fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a1_a_aq,fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({vcc,vcc,vcc}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.ax_width = 22;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.ay_scan_in_width = 15;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.operation_mode = "m27x27";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.result_a_width = 37;
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.signed_max = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "90A736506F4DD878815EDA844CDDF7B62798C2CEDD2A0C6A82D26AF452A470BF";

fourteennm_lcell_comb fp_functions_0_aadd_11_a122(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_11_a127_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_11_a122_cout),
	.shareout());
defparam fp_functions_0_aadd_11_a122.extended_lut = "off";
defparam fp_functions_0_aadd_11_a122.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a122.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a37.extended_lut = "off";
defparam fp_functions_0_aadd_2_a37.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a37.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai112_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai116_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai116_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai116_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "2ACF76DAEC62BF463B51BF0690852D1EC74F5BF80C55865FAFC52669990BDA68";

fourteennm_lcell_comb fp_functions_0_aadd_11_a127(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_11_a127_cout),
	.shareout());
defparam fp_functions_0_aadd_11_a127.extended_lut = "off";
defparam fp_functions_0_aadd_11_a127.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_11_a127.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a42.extended_lut = "off";
defparam fp_functions_0_aadd_2_a42.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_2_a42.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_lowRangeB_uid74_invPolyEval_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_lowRangeB_uid74_invPolyEval_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist5_lowRangeB_uid74_invPolyEval_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_lowRangeB_uid74_invPolyEval_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a0_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a1_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a2_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a3_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a4_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a5_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a6_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a7_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a8_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a9_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a10_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a11_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a12_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a13_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a14_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a15_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a16_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a17_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a18_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a19_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a20_a_aq));
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a8_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a9_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a10_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a11_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a12_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a13_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a14_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a14_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1326_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist1_yaddr_uid36_fpinversetest_merged_bit_select_b_14_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ram_block fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC0_uid60_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC0_uid60_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 29;
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC0_uid60_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "0C9C9C3A0E08374926D19F5D595A68D1C5A0EA5B4846A61A10053FB1EB7F34E0";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a47.extended_lut = "off";
defparam fp_functions_0_aadd_2_a47.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_2_a47.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_6_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a1_sumout),
	.cout(fp_functions_0_aadd_6_a2),
	.shareout());
defparam fp_functions_0_aadd_6_a1.extended_lut = "off";
defparam fp_functions_0_aadd_6_a1.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a6_sumout),
	.cout(fp_functions_0_aadd_6_a7),
	.shareout());
defparam fp_functions_0_aadd_6_a6.extended_lut = "off";
defparam fp_functions_0_aadd_6_a6.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a11_sumout),
	.cout(fp_functions_0_aadd_6_a12),
	.shareout());
defparam fp_functions_0_aadd_6_a11.extended_lut = "off";
defparam fp_functions_0_aadd_6_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a16_sumout),
	.cout(fp_functions_0_aadd_6_a17),
	.shareout());
defparam fp_functions_0_aadd_6_a16.extended_lut = "off";
defparam fp_functions_0_aadd_6_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a21_sumout),
	.cout(fp_functions_0_aadd_6_a22),
	.shareout());
defparam fp_functions_0_aadd_6_a21.extended_lut = "off";
defparam fp_functions_0_aadd_6_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a26_sumout),
	.cout(fp_functions_0_aadd_6_a27),
	.shareout());
defparam fp_functions_0_aadd_6_a26.extended_lut = "off";
defparam fp_functions_0_aadd_6_a26.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a31_sumout),
	.cout(fp_functions_0_aadd_6_a32),
	.shareout());
defparam fp_functions_0_aadd_6_a31.extended_lut = "off";
defparam fp_functions_0_aadd_6_a31.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a36_sumout),
	.cout(fp_functions_0_aadd_6_a37),
	.shareout());
defparam fp_functions_0_aadd_6_a36.extended_lut = "off";
defparam fp_functions_0_aadd_6_a36.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a41_sumout),
	.cout(fp_functions_0_aadd_6_a42),
	.shareout());
defparam fp_functions_0_aadd_6_a41.extended_lut = "off";
defparam fp_functions_0_aadd_6_a41.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a46_sumout),
	.cout(fp_functions_0_aadd_6_a47),
	.shareout());
defparam fp_functions_0_aadd_6_a46.extended_lut = "off";
defparam fp_functions_0_aadd_6_a46.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a51_sumout),
	.cout(fp_functions_0_aadd_6_a52),
	.shareout());
defparam fp_functions_0_aadd_6_a51.extended_lut = "off";
defparam fp_functions_0_aadd_6_a51.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a56_sumout),
	.cout(fp_functions_0_aadd_6_a57),
	.shareout());
defparam fp_functions_0_aadd_6_a56.extended_lut = "off";
defparam fp_functions_0_aadd_6_a56.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a61(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a61_sumout),
	.cout(fp_functions_0_aadd_6_a62),
	.shareout());
defparam fp_functions_0_aadd_6_a61.extended_lut = "off";
defparam fp_functions_0_aadd_6_a61.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a66(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a66_sumout),
	.cout(fp_functions_0_aadd_6_a67),
	.shareout());
defparam fp_functions_0_aadd_6_a66.extended_lut = "off";
defparam fp_functions_0_aadd_6_a66.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a71(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a71_sumout),
	.cout(fp_functions_0_aadd_6_a72),
	.shareout());
defparam fp_functions_0_aadd_6_a71.extended_lut = "off";
defparam fp_functions_0_aadd_6_a71.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a76(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a76_sumout),
	.cout(fp_functions_0_aadd_6_a77),
	.shareout());
defparam fp_functions_0_aadd_6_a76.extended_lut = "off";
defparam fp_functions_0_aadd_6_a76.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a81(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a81_sumout),
	.cout(fp_functions_0_aadd_6_a82),
	.shareout());
defparam fp_functions_0_aadd_6_a81.extended_lut = "off";
defparam fp_functions_0_aadd_6_a81.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a86(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a86_sumout),
	.cout(fp_functions_0_aadd_6_a87),
	.shareout());
defparam fp_functions_0_aadd_6_a86.extended_lut = "off";
defparam fp_functions_0_aadd_6_a86.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a91(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a91_sumout),
	.cout(fp_functions_0_aadd_6_a92),
	.shareout());
defparam fp_functions_0_aadd_6_a91.extended_lut = "off";
defparam fp_functions_0_aadd_6_a91.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a96(
	.dataa(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a96_sumout),
	.cout(fp_functions_0_aadd_6_a97),
	.shareout());
defparam fp_functions_0_aadd_6_a96.extended_lut = "off";
defparam fp_functions_0_aadd_6_a96.lut_mask = 64'h00000000005555AA;
defparam fp_functions_0_aadd_6_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a101_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_6_a101.extended_lut = "off";
defparam fp_functions_0_aadd_6_a101.lut_mask = 64'h0000000000000FF0;
defparam fp_functions_0_aadd_6_a101.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_mac fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a11_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a10_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a9_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a8_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a7_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a6_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a5_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a4_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a3_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a2_a_aq,fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a1_a_aq,
fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({areset,areset}),
	.ena({vcc,vcc,vcc}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.ax_width = 12;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.ay_scan_in_width = 12;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.az_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.by_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.operation_mode = "m18x18_full";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.output_clock = "1";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.result_a_width = 24;
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.signed_max = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.signed_may = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "EE11525F7D0F5E66F88981669C3C1AFDE4D22085EE6809A5A9F66C3154CDA6BA";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "0D6EEF2B5B7EC8FD9AC5B7E904E608D01523AF869EC6F48B79FC66A5B7093336";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "03E435912296FC120FBED22F549D3F08BC7261E787D34EBC51283C171773F885";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "5D0C843CA1C54B1237A4772957B033214A356F1057CEC0E16C7C86F8BD093C32";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "6B09868162B932E62F19E06C89AED2DC48D40394FE585952EDC7BCF5265984A8";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "725B872B1CD4FCAE357EAFBBEBB5E6146749083610D72912551B5BC05E0AE02E";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "7C6D2D6700E6AA61C6559FCD5846AE19206B0D774F7059B338E8421110E5DB42";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "7F8E364A55AD99E007992AA4C7F8CB4B1F8DA4F795306C8C540D3CB1B0A142F6";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "7FF038739936D2B552B4999C3FFF0C6DAAA49C0819A5247F995B00DB70CB3CAE";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "D5556AD6B4924993318C787C00000F8E3336D6AAB4931C001E6DAA48F0F2559E";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "9999B364D92492DA5AD6AD56AAAAA55A96924D998C70FC001F8E336D5A56CC7E";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "E1E1C3871E38E31C6318CE673333366CDB2496D2D6A556AAB55A96DB3631C3FE";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "FE01FC07E03F03E07C1F0F87C3C3C78F1C38E71CE73998CCD99324925B5A9554";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "FFFE0007FFC003FF801FF007FC03F80FE03F07E0F83E1F0F1E1C38E39C631998";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "FFFFFFF8000003FFFFE00007FFFC000FFFC007FF003FE00FE01FC0FC1F83E1E0";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "FFFFFFFFFFFFFC0000000007FFFFFFF0000007FFFFC0000FFFE000FFE003FE00";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFF800000000000007FFFFFFFFF0000000FFFFFC0000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "00000000000000000000000000000000000007FFFFFFFFFFFFFFFF0000000000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000";

fourteennm_ram_block fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC1_uid63_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fp_functions_0|memoryC1_uid63_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 20;
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC1_uid63_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1063_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 3;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 4;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 5;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fp_functions_0|redist3_yaddr_uid36_fpinversetest_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 15;
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1334_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1334_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1334_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a7_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a0_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a1_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a2_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a3_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a4_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a5_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a6_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a7_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a8_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a9_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a10_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a11_a_aq));
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1071_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1071_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1071_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a0_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a1_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a2_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a2_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai825_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fp_functions_0|redist0_yaddr_uid36_fpinversetest_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a8_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "A4C38078760372CB4DB0518569CB0244C3A2AFF74309ECD2F7718E4A5A84DC0C";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "9E57B2E6BD265E53D0ADC629857BBD947469E351DEF10D69B0AEFFD9A8C320E2";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "FDCF6E118F113649349BD284ABD112A1594D2B9DE2F9EC380B6A2971D7CE828F";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "83C0E1F07CF0F1C70C78CE6398C8899334DB794B57ACB952D24CCE7E003E665A";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "803FE00FFC0FF03F03F83E1F87C7878F0C38E738CE6464C9B6DA5AD55554B493";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "80001FFFFC000FFF0007FE007FC07F80FC07E0F83E1C1C3871C639CCCCCD9249";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "8000000003FFFFFF000001FFFFC0007FFC001FF801FC03F80FC1F83C3C3C71C7";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "8000000000000000FFFFFFFFFFC0000003FFFFF80003FFF8003FF803FC03F03F";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "7FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000007FFFFFFF8000007FFFC000FFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "000000000000000000000000003FFFFFFFFFFFFFFFFFFFF80000000003FFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFF";

fourteennm_ram_block fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(gnd),
	.aclr(gnd),
	.sclr(areset),
	.ena0(vcc),
	.ena1(vcc),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15]}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fp_functions_191/synth/Float_Inv_altera_fp_functions_191_j4yadhq_memoryC2_uid66_inverseTables_lutmem.hex";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fp_functions_0|memoryC2_uid66_inverseTables_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock0";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 12;
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fp_functions_0_amemoryC2_uid66_inverseTables_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a3_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a4_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a5_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a6_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a7_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a8_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a9_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a10_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a11_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a12_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a13_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a14_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a0_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a1_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a2_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_1_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a9_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a3_a(
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a3_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a4_a(
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a4_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a5_a(
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a5_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a6_a(
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a6_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a7_a(
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a7_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a8_a(
	.clk(clk),
	.d(a[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a8_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a9_a(
	.clk(clk),
	.d(a[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a9_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a10_a(
	.clk(clk),
	.d(a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a10_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a11_a(
	.clk(clk),
	.d(a[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a11_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a12_a(
	.clk(clk),
	.d(a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a12_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a13_a(
	.clk(clk),
	.d(a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a13_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a14_a(
	.clk(clk),
	.d(a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a14_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a0_a(
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a0_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a1_a(
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a1_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a2_a(
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a2_a_aq));
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_delay_0_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai833_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai833_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai833_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a10_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a11_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a12_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a13_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid23_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a14_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a15_a_a0_a_aq));
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aMux_32_a2(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a0_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_32_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_32_a2.extended_lut = "off";
defparam fp_functions_0_aMux_32_a2.lut_mask = 64'h4000D57F4000D57F;
defparam fp_functions_0_aMux_32_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_31_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_31_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_31_a0.extended_lut = "off";
defparam fp_functions_0_aMux_31_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_31_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_30_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a2_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_30_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_30_a0.extended_lut = "off";
defparam fp_functions_0_aMux_30_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_30_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_29_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a3_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_29_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_29_a0.extended_lut = "off";
defparam fp_functions_0_aMux_29_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_29_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_28_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_28_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_28_a0.extended_lut = "off";
defparam fp_functions_0_aMux_28_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_28_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_27_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a5_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_27_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_27_a0.extended_lut = "off";
defparam fp_functions_0_aMux_27_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_27_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_26_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_26_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_26_a0.extended_lut = "off";
defparam fp_functions_0_aMux_26_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_26_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_25_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a7_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_25_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_25_a0.extended_lut = "off";
defparam fp_functions_0_aMux_25_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_25_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_24_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a8_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_24_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_24_a0.extended_lut = "off";
defparam fp_functions_0_aMux_24_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_24_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_23_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a9_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_23_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_23_a0.extended_lut = "off";
defparam fp_functions_0_aMux_23_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_23_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_22_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a10_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_22_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_22_a0.extended_lut = "off";
defparam fp_functions_0_aMux_22_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_22_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_21_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a11_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_21_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_21_a0.extended_lut = "off";
defparam fp_functions_0_aMux_21_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_21_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_20_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a12_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_20_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_20_a0.extended_lut = "off";
defparam fp_functions_0_aMux_20_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_20_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_19_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a13_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_19_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_19_a0.extended_lut = "off";
defparam fp_functions_0_aMux_19_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_19_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_18_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a14_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_18_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_18_a0.extended_lut = "off";
defparam fp_functions_0_aMux_18_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_18_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_17_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a15_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_17_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_17_a0.extended_lut = "off";
defparam fp_functions_0_aMux_17_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_17_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_16_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a16_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_16_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_16_a0.extended_lut = "off";
defparam fp_functions_0_aMux_16_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_16_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_15_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a17_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_15_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_15_a0.extended_lut = "off";
defparam fp_functions_0_aMux_15_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_15_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_14_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a18_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_14_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_14_a0.extended_lut = "off";
defparam fp_functions_0_aMux_14_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_14_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_13_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a19_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_13_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_13_a0.extended_lut = "off";
defparam fp_functions_0_aMux_13_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_13_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_12_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a20_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_12_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_12_a0.extended_lut = "off";
defparam fp_functions_0_aMux_12_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_12_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_11_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a21_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_11_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_11_a0.extended_lut = "off";
defparam fp_functions_0_aMux_11_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_11_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_10_a0(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a22_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_10_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_10_a0.extended_lut = "off";
defparam fp_functions_0_aMux_10_a0.lut_mask = 64'h0000957F0000957F;
defparam fp_functions_0_aMux_10_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a2(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a0_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a2.extended_lut = "off";
defparam fp_functions_0_aMux_9_a2.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a3(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a3.extended_lut = "off";
defparam fp_functions_0_aMux_9_a3.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a4(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a2_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a4.extended_lut = "off";
defparam fp_functions_0_aMux_9_a4.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a5(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a3_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a5.extended_lut = "off";
defparam fp_functions_0_aMux_9_a5.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a6(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a6.extended_lut = "off";
defparam fp_functions_0_aMux_9_a6.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a7(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a5_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a7.extended_lut = "off";
defparam fp_functions_0_aMux_9_a7.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a8(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a6_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a8.extended_lut = "off";
defparam fp_functions_0_aMux_9_a8.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_9_a9(
	.dataa(!fp_functions_0_aredist7_excN_x_uid26_fpInverseTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aexcI_x_uid25_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fp_functions_0_axRegAndUdf_uid49_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aredist9_excZ_x_uid21_fpInverseTest_q_1_q_a0_a_aq),
	.datae(!fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_o_a7_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_9_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_9_a9.extended_lut = "off";
defparam fp_functions_0_aMux_9_a9.lut_mask = 64'h4080D5FF4080D5FF;
defparam fp_functions_0_aMux_9_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_3_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datae(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_3_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_3_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_3_a0.lut_mask = 64'h0000000100000001;
defparam fp_functions_0_areduce_nor_3_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(!fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a.lut_mask = 64'h0000010000000100;
defparam fp_functions_0_aexcN_x_uid26_fpInverseTest_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(!fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a.lut_mask = 64'h0000000100000001;
defparam fp_functions_0_aexcI_x_uid25_fpInverseTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_5_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.datae(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_5_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_5_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_5_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_5_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_a0_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(!fp_functions_0_aadd_2_a1_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0.lut_mask = 64'h00000000FFFE7F7E;
defparam fp_functions_0_axRegAndUdf_uid49_fpInverseTest_qi_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_5(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_5_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_5.extended_lut = "off";
defparam fp_functions_0_areduce_nor_5.lut_mask = 64'h0080008000800080;
defparam fp_functions_0_areduce_nor_5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0.extended_lut = "off";
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_afracRCalc_uid47_fpInverseTest_q_a6_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.datad(!fp_functions_0_aredist8_fracXIsZero_uid23_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datae(!fp_functions_0_aredist10_singX_uid8_fpInverseTest_b_16_adelay_signals_a0_a_a0_a_aq),
	.dataf(!fp_functions_0_areduce_nor_3_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a.lut_mask = 64'h0000FFFF0000FEFF;
defparam fp_functions_0_asignR_uid57_fpInverseTest_qi_a0_a.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a36_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.datab(!fp_functions_0_aredist6_fracXIsZero_uid31_fpInverseTest_q_16_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0.extended_lut = "off";
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_aexpRCompYIsOneExt_uid42_fpInverseTest_expRCalc_uid48_fpInverseTest_merged_a1_a1_a_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai138_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai138_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai138_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_wraddr_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(a[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai100_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai102_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_sticky_ena_q_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_cmpReg_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai102_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai102_a0.extended_lut = "off";
defparam fp_functions_0_ai102_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai102_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(a[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(a[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(a[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(a[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(a[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(a[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(a[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai138_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai138_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai138_a0.extended_lut = "off";
defparam fp_functions_0_ai138_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai138_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai138_a1(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai138_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai138_a1.extended_lut = "off";
defparam fp_functions_0_ai138_a1.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai138_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai138_a2(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai138_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai138_a2.extended_lut = "off";
defparam fp_functions_0_ai138_a2.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai138_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai100_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq),
	.datae(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai100_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai100_a0.extended_lut = "off";
defparam fp_functions_0_ai100_a0.lut_mask = 64'h0000002000000020;
defparam fp_functions_0_ai100_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist5_lowRangeB_uid74_invPolyEval_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_as1sumAHighB_uid76_invPolyEval_o_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ch_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_ai100_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq_aq));
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai112_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai112_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai112_a0.extended_lut = "off";
defparam fp_functions_0_ai112_a0.lut_mask = 64'h9999999999999999;
defparam fp_functions_0_ai112_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai116_a0(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai116_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai116_a0.extended_lut = "off";
defparam fp_functions_0_ai116_a0.lut_mask = 64'h6C6C6C6C6C6C6C6C;
defparam fp_functions_0_ai116_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai116_a1(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai116_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai116_a1.extended_lut = "off";
defparam fp_functions_0_ai116_a1.lut_mask = 64'h1E3C1E3C1E3C1E3C;
defparam fp_functions_0_ai116_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai116_a2(
	.dataa(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_i_a3_a_aq),
	.datae(!fp_functions_0_aredist11_expX_uid6_fpInverseTest_b_16_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai116_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai116_a2.extended_lut = "off";
defparam fp_functions_0_ai116_a2.lut_mask = 64'h01FE03FC01FE03FC;
defparam fp_functions_0_ai116_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid88_pT2_uid79_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1348_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1324_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1326_a0(
	.dataa(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_sticky_ena_q_a0_a_aq),
	.datab(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_cmpReg_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1326_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1326_a0.extended_lut = "off";
defparam fp_functions_0_ai1326_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai1326_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1348_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1348_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1348_a0.extended_lut = "off";
defparam fp_functions_0_ai1348_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai1348_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1324_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1324_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1324_a0.extended_lut = "off";
defparam fp_functions_0_ai1324_a0.lut_mask = 64'h0200020002000200;
defparam fp_functions_0_ai1324_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_memoryC2_uid66_inverseTables_lutmem_r_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aprodXY_uid85_pT1_uid73_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1085_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1061_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1063_a0(
	.dataa(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.datab(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_cmpReg_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1063_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1063_a0.extended_lut = "off";
defparam fp_functions_0_ai1063_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai1063_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist2_yAddr_uid36_fpInverseTest_merged_bit_select_c_3_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_ai1324_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq_aq));
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1334_a0(
	.dataa(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1334_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1334_a0.extended_lut = "off";
defparam fp_functions_0_ai1334_a0.lut_mask = 64'h9999999999999999;
defparam fp_functions_0_ai1334_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1334_a1(
	.dataa(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1334_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1334_a1.extended_lut = "off";
defparam fp_functions_0_ai1334_a1.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai1334_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1334_a2(
	.dataa(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist1_yAddr_uid36_fpInverseTest_merged_bit_select_b_14_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1334_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1334_a2.extended_lut = "off";
defparam fp_functions_0_ai1334_a2.lut_mask = 64'h1EF01EF01EF01EF0;
defparam fp_functions_0_ai1334_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1085_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1085_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1085_a0.extended_lut = "off";
defparam fp_functions_0_ai1085_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai1085_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1061_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1061_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1061_a0.extended_lut = "off";
defparam fp_functions_0_ai1061_a0.lut_mask = 64'h0200020002000200;
defparam fp_functions_0_ai1061_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_ai1061_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq_aq));
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1071_a0(
	.dataa(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1071_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1071_a0.extended_lut = "off";
defparam fp_functions_0_ai1071_a0.lut_mask = 64'h9999999999999999;
defparam fp_functions_0_ai1071_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1071_a1(
	.dataa(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1071_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1071_a1.extended_lut = "off";
defparam fp_functions_0_ai1071_a1.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai1071_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1071_a2(
	.dataa(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist3_yAddr_uid36_fpInverseTest_merged_bit_select_c_10_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1071_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1071_a2.extended_lut = "off";
defparam fp_functions_0_ai1071_a2.lut_mask = 64'h1EF01EF01EF01EF0;
defparam fp_functions_0_ai1071_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai847_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_cmpReg_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai823_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_cmpReg_q_a0_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai825_a0(
	.dataa(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_cmpReg_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai825_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai825_a0.extended_lut = "off";
defparam fp_functions_0_ai825_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai825_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(a[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(a[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(a[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai847_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai847_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai847_a0.extended_lut = "off";
defparam fp_functions_0_ai847_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_ai847_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai823_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datac(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datad(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai823_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai823_a0.extended_lut = "off";
defparam fp_functions_0_ai823_a0.lut_mask = 64'h0200020002000200;
defparam fp_functions_0_ai823_a0.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq(
	.clk(clk),
	.d(fp_functions_0_ai823_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq_aq));
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai833_a0(
	.dataa(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai833_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai833_a0.extended_lut = "off";
defparam fp_functions_0_ai833_a0.lut_mask = 64'h9999999999999999;
defparam fp_functions_0_ai833_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai833_a1(
	.dataa(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai833_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai833_a1.extended_lut = "off";
defparam fp_functions_0_ai833_a1.lut_mask = 64'h6363636363636363;
defparam fp_functions_0_ai833_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai833_a2(
	.dataa(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datab(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datac(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datad(!fp_functions_0_aredist0_yAddr_uid36_fpInverseTest_merged_bit_select_b_7_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai833_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai833_a2.extended_lut = "off";
defparam fp_functions_0_ai833_a2.lut_mask = 64'h1EF01EF01EF01EF0;
defparam fp_functions_0_ai833_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_afracXIsZero_uid23_fpInverseTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid23_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid23_fpInverseTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid23_fpInverseTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0(
	.dataa(!areset),
	.datab(!a[3]),
	.datac(!a[0]),
	.datad(!a[1]),
	.datae(!a[2]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0.extended_lut = "off";
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1(
	.dataa(!a[5]),
	.datab(!a[6]),
	.datac(!a[7]),
	.datad(!a[8]),
	.datae(!a[9]),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1.extended_lut = "off";
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2(
	.dataa(!a[15]),
	.datab(!a[16]),
	.datac(!a[11]),
	.datad(!a[12]),
	.datae(!a[13]),
	.dataf(!a[14]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2.extended_lut = "off";
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3(
	.dataa(!a[17]),
	.datab(!a[18]),
	.datac(!a[19]),
	.datad(!a[20]),
	.datae(!a[21]),
	.dataf(!a[22]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3.extended_lut = "off";
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4(
	.dataa(!a[4]),
	.datab(!a[10]),
	.datac(!fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a0_combout),
	.datad(!fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a1_combout),
	.datae(!fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a2_combout),
	.dataf(!fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4.extended_lut = "off";
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4.lut_mask = 64'h0000000000000008;
defparam fp_functions_0_afracXIsZero_uid31_fpInverseTest_delay_ai6_a4.shared_arith = "off";

assign q[22] = fp_functions_0_aMux_10_a0_combout;

assign q[21] = fp_functions_0_aMux_11_a0_combout;

assign q[20] = fp_functions_0_aMux_12_a0_combout;

assign q[19] = fp_functions_0_aMux_13_a0_combout;

assign q[18] = fp_functions_0_aMux_14_a0_combout;

assign q[17] = fp_functions_0_aMux_15_a0_combout;

assign q[16] = fp_functions_0_aMux_16_a0_combout;

assign q[15] = fp_functions_0_aMux_17_a0_combout;

assign q[14] = fp_functions_0_aMux_18_a0_combout;

assign q[13] = fp_functions_0_aMux_19_a0_combout;

assign q[12] = fp_functions_0_aMux_20_a0_combout;

assign q[11] = fp_functions_0_aMux_21_a0_combout;

assign q[10] = fp_functions_0_aMux_22_a0_combout;

assign q[9] = fp_functions_0_aMux_23_a0_combout;

assign q[8] = fp_functions_0_aMux_24_a0_combout;

assign q[7] = fp_functions_0_aMux_25_a0_combout;

assign q[6] = fp_functions_0_aMux_26_a0_combout;

assign q[5] = fp_functions_0_aMux_27_a0_combout;

assign q[4] = fp_functions_0_aMux_28_a0_combout;

assign q[3] = fp_functions_0_aMux_29_a0_combout;

assign q[2] = fp_functions_0_aMux_30_a0_combout;

assign q[1] = fp_functions_0_aMux_31_a0_combout;

assign q[0] = fp_functions_0_aMux_32_a2_combout;

assign q[23] = fp_functions_0_aMux_9_a2_combout;

assign q[24] = fp_functions_0_aMux_9_a3_combout;

assign q[25] = fp_functions_0_aMux_9_a4_combout;

assign q[26] = fp_functions_0_aMux_9_a5_combout;

assign q[27] = fp_functions_0_aMux_9_a6_combout;

assign q[28] = fp_functions_0_aMux_9_a7_combout;

assign q[29] = fp_functions_0_aMux_9_a8_combout;

assign q[30] = fp_functions_0_aMux_9_a9_combout;

assign q[31] = fp_functions_0_asignR_uid57_fpInverseTest_delay_adelay_signals_a0_a_a0_a_aq;

endmodule
