// Float_MulAdd.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module Float_MulAdd (
		input  wire        clk,    //    clk.clk
		input  wire        areset, // areset.reset
		input  wire [31:0] a,      //      a.a
		input  wire [31:0] b,      //      b.b
		input  wire [31:0] c,      //      c.c
		output wire [31:0] q       //      q.q
	);

	Float_MulAdd_altera_fp_functions_191_e2g3mei fp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.areset (areset), //   input,   width = 1, areset.reset
		.a      (a),      //   input,  width = 32,      a.a
		.b      (b),      //   input,  width = 32,      b.b
		.c      (c),      //   input,  width = 32,      c.c
		.q      (q)       //  output,  width = 32,      q.q
	);

endmodule
