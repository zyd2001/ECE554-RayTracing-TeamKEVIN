module IC_Controller();

endmodule