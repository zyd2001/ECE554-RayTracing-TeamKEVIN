// Fix_Div.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module Fix_Div (
		input  wire        clk,         //         clk.clk
		input  wire        rst,         //         rst.reset
		input  wire [0:0]  en,          //          en.en
		input  wire [31:0] numerator,   //   numerator.numerator
		input  wire [31:0] denominator, // denominator.denominator
		output wire [31:0] result       //      result.result
	);

	Fix_Div_altera_fxp_functions_191_fy4uury fxp_functions_0 (
		.clk         (clk),         //   input,   width = 1,         clk.clk
		.rst         (rst),         //   input,   width = 1,         rst.reset
		.en          (en),          //   input,   width = 1,          en.en
		.numerator   (numerator),   //   input,  width = 32,   numerator.numerator
		.denominator (denominator), //   input,  width = 32, denominator.denominator
		.result      (result)       //  output,  width = 32,      result.result
	);

endmodule
