// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/20/2021 23:00:20"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module ItoF (
	q,
	clk,
	areset,
	en,
	a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	clk;
input 	areset;
input 	[0:0] en;
input 	[31:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a0_a_aq;
wire fp_functions_0_aadd_4_a1_sumout;
wire fp_functions_0_aadd_5_a1_sumout;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a8_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a9_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a10_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a11_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a12_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a13_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a14_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a15_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a16_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a17_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a18_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a19_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a20_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a21_a_aq;
wire fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a22_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_ainIsZero_uid12_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aadd_3_a1_sumout;
wire fp_functions_0_aadd_3_a2;
wire fp_functions_0_aadd_4_a7_cout;
wire fp_functions_0_aadd_5_a7_cout;
wire fp_functions_0_aadd_3_a6_sumout;
wire fp_functions_0_aadd_3_a7;
wire fp_functions_0_aadd_3_a11_sumout;
wire fp_functions_0_aadd_3_a12;
wire fp_functions_0_aadd_3_a16_sumout;
wire fp_functions_0_aadd_3_a17;
wire fp_functions_0_aadd_3_a21_sumout;
wire fp_functions_0_aadd_3_a22;
wire fp_functions_0_aadd_3_a26_sumout;
wire fp_functions_0_aadd_3_a27;
wire fp_functions_0_aadd_3_a31_sumout;
wire fp_functions_0_aadd_3_a32;
wire fp_functions_0_aadd_3_a36_sumout;
wire fp_functions_0_aadd_3_a37;
wire fp_functions_0_aadd_3_a41_sumout;
wire fp_functions_0_aadd_3_a42;
wire fp_functions_0_aadd_3_a46_sumout;
wire fp_functions_0_aadd_3_a47;
wire fp_functions_0_aadd_3_a51_sumout;
wire fp_functions_0_aadd_3_a52;
wire fp_functions_0_aadd_3_a56_sumout;
wire fp_functions_0_aadd_3_a57;
wire fp_functions_0_aadd_3_a61_sumout;
wire fp_functions_0_aadd_3_a62;
wire fp_functions_0_aadd_3_a66_sumout;
wire fp_functions_0_aadd_3_a67;
wire fp_functions_0_aadd_3_a71_sumout;
wire fp_functions_0_aadd_3_a72;
wire fp_functions_0_aadd_3_a76_sumout;
wire fp_functions_0_aadd_3_a77;
wire fp_functions_0_aadd_3_a81_sumout;
wire fp_functions_0_aadd_3_a82;
wire fp_functions_0_aadd_3_a86_sumout;
wire fp_functions_0_aadd_3_a87;
wire fp_functions_0_aadd_3_a91_sumout;
wire fp_functions_0_aadd_3_a92;
wire fp_functions_0_aadd_3_a96_sumout;
wire fp_functions_0_aadd_3_a97;
wire fp_functions_0_aadd_3_a101_sumout;
wire fp_functions_0_aadd_3_a102;
wire fp_functions_0_aadd_3_a106_sumout;
wire fp_functions_0_aadd_3_a107;
wire fp_functions_0_aadd_3_a111_sumout;
wire fp_functions_0_aadd_3_a112;
wire fp_functions_0_aadd_3_a116_sumout;
wire fp_functions_0_aadd_3_a117;
wire fp_functions_0_aadd_3_a121_sumout;
wire fp_functions_0_aadd_3_a122;
wire fp_functions_0_aadd_3_a126_sumout;
wire fp_functions_0_aadd_3_a127;
wire fp_functions_0_aadd_3_a131_sumout;
wire fp_functions_0_aadd_3_a132;
wire fp_functions_0_aadd_3_a136_sumout;
wire fp_functions_0_aadd_3_a137;
wire fp_functions_0_aadd_3_a141_sumout;
wire fp_functions_0_aadd_3_a142;
wire fp_functions_0_aadd_3_a146_sumout;
wire fp_functions_0_aadd_3_a147;
wire fp_functions_0_aadd_3_a151_sumout;
wire fp_functions_0_aadd_3_a152;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a1_a_a0_a_aq;
wire fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a_aq;
wire fp_functions_0_aadd_3_a157_cout;
wire fp_functions_0_aadd_4_a12_cout;
wire fp_functions_0_aadd_5_a12_cout;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a2_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a3_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a4_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a5_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a6_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a7_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a8_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a9_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a10_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a11_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a12_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a13_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a14_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a15_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a16_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a17_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a18_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a19_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a20_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a21_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a22_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a23_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a0_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a1_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a2_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a3_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a4_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a5_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a6_a_aq;
wire fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a7_a_aq;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a2_a_a0_a_aq;
wire fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_1_a0_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq;
wire fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a_aq;
wire fp_functions_0_asticky_uid20_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a_aq;
wire fp_functions_0_aadd_4_a17_cout;
wire fp_functions_0_aadd_5_a17_cout;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq;
wire fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq;
wire fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq;
wire fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a_aq;
wire fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a_aq;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a3_a_a0_a_aq;
wire fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_0_a0_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq;
wire fp_functions_0_aadd_3_a161_sumout;
wire fp_functions_0_aadd_4_a22_cout;
wire fp_functions_0_aadd_5_a22_cout;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq;
wire fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_aq;
wire fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_1_a0_a_aq;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a4_a_a0_a_aq;
wire fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq;
wire fp_functions_0_aadd_4_a27_cout;
wire fp_functions_0_aadd_5_a27_cout;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq;
wire fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_0_a0_a_aq;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a5_a_a0_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a_aq;
wire fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a_aq;
wire fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a_aq;
wire fp_functions_0_aadd_4_a32_cout;
wire fp_functions_0_aadd_5_a32_cout;
wire fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a6_a_a0_a_aq;
wire fp_functions_0_aadd_0_a1_sumout;
wire fp_functions_0_aadd_0_a2;
wire fp_functions_0_aadd_0_a6_sumout;
wire fp_functions_0_aadd_0_a7;
wire fp_functions_0_aadd_0_a11_sumout;
wire fp_functions_0_aadd_0_a12;
wire fp_functions_0_aadd_0_a16_sumout;
wire fp_functions_0_aadd_0_a17;
wire fp_functions_0_aadd_0_a21_sumout;
wire fp_functions_0_aadd_0_a22;
wire fp_functions_0_aadd_0_a26_sumout;
wire fp_functions_0_aadd_0_a27;
wire fp_functions_0_aadd_0_a31_sumout;
wire fp_functions_0_aadd_0_a32;
wire fp_functions_0_aadd_0_a36_sumout;
wire fp_functions_0_aadd_0_a37;
wire fp_functions_0_aadd_0_a41_sumout;
wire fp_functions_0_aadd_0_a42;
wire fp_functions_0_aadd_0_a46_sumout;
wire fp_functions_0_aadd_0_a47;
wire fp_functions_0_aadd_0_a51_sumout;
wire fp_functions_0_aadd_0_a52;
wire fp_functions_0_aadd_0_a56_sumout;
wire fp_functions_0_aadd_0_a57;
wire fp_functions_0_aadd_0_a61_sumout;
wire fp_functions_0_aadd_0_a62;
wire fp_functions_0_aadd_0_a66_sumout;
wire fp_functions_0_aadd_0_a67;
wire fp_functions_0_aadd_0_a71_sumout;
wire fp_functions_0_aadd_0_a72;
wire fp_functions_0_aadd_0_a76_sumout;
wire fp_functions_0_aadd_0_a77;
wire fp_functions_0_aadd_0_a81_sumout;
wire fp_functions_0_aadd_0_a82;
wire fp_functions_0_aadd_0_a86_sumout;
wire fp_functions_0_aadd_0_a87;
wire fp_functions_0_aadd_0_a91_sumout;
wire fp_functions_0_aadd_0_a92;
wire fp_functions_0_aadd_0_a96_sumout;
wire fp_functions_0_aadd_0_a97;
wire fp_functions_0_aadd_0_a101_sumout;
wire fp_functions_0_aadd_0_a102;
wire fp_functions_0_aadd_0_a106_sumout;
wire fp_functions_0_aadd_0_a107;
wire fp_functions_0_aadd_0_a111_sumout;
wire fp_functions_0_aadd_0_a112;
wire fp_functions_0_aadd_0_a116_sumout;
wire fp_functions_0_aadd_0_a117;
wire fp_functions_0_aadd_0_a121_sumout;
wire fp_functions_0_aadd_0_a122;
wire fp_functions_0_aadd_0_a126_sumout;
wire fp_functions_0_aadd_0_a127;
wire fp_functions_0_aadd_0_a131_sumout;
wire fp_functions_0_aadd_0_a132;
wire fp_functions_0_aadd_0_a136_sumout;
wire fp_functions_0_aadd_0_a141_sumout;
wire fp_functions_0_aadd_0_a142;
wire fp_functions_0_aadd_0_a146_sumout;
wire fp_functions_0_aadd_0_a147;
wire fp_functions_0_aadd_0_a151_sumout;
wire fp_functions_0_aadd_0_a152;
wire fp_functions_0_aadd_0_a156_sumout;
wire fp_functions_0_aadd_0_a157;
wire fp_functions_0_aadd_4_a37_cout;
wire fp_functions_0_aadd_5_a37_cout;
wire fp_functions_0_aadd_4_a42_cout;
wire fp_functions_0_aadd_5_a42_cout;
wire fp_functions_0_aadd_4_a47_cout;
wire fp_functions_0_aadd_5_a47_cout;
wire fp_functions_0_ai1302_a10_cout;
wire fp_functions_0_ai1302_a14_sumout;
wire fp_functions_0_ai1302_a15;
wire fp_functions_0_ai1302_a19_sumout;
wire fp_functions_0_ai1302_a20;
wire fp_functions_0_ai1302_a24_sumout;
wire fp_functions_0_ai1302_a25;
wire fp_functions_0_ai1302_a29_sumout;
wire fp_functions_0_ai1302_a30;
wire fp_functions_0_ai1302_a34_sumout;
wire fp_functions_0_ai1302_a35;
wire fp_functions_0_ai1302_a39_sumout;
wire fp_functions_0_ai1302_a40;
wire fp_functions_0_ai1302_a44_sumout;
wire fp_functions_0_ai1302_a45;
wire fp_functions_0_ai1302_a49_sumout;
wire fp_functions_0_ai1302_a50;
wire fp_functions_0_ai1302_a54_sumout;
wire fp_functions_0_ai1302_a55;
wire fp_functions_0_ai1302_a59_sumout;
wire fp_functions_0_ai1302_a60;
wire fp_functions_0_ai1302_a64_sumout;
wire fp_functions_0_ai1302_a70_cout;
wire fp_functions_0_ai1302_a74_sumout;
wire fp_functions_0_ai1302_a75;
wire fp_functions_0_ai1302_a79_sumout;
wire fp_functions_0_ai1302_a80;
wire fp_functions_0_ai1302_a84_sumout;
wire fp_functions_0_ai1302_a85;
wire fp_functions_0_ai1302_a89_sumout;
wire fp_functions_0_ai1302_a90;
wire fp_functions_0_ai1302_a94_sumout;
wire fp_functions_0_ai1302_a95;
wire fp_functions_0_ai1302_a99_sumout;
wire fp_functions_0_ai1302_a100;
wire fp_functions_0_ai1302_a104_sumout;
wire fp_functions_0_ai1302_a105;
wire fp_functions_0_ai1302_a109_sumout;
wire fp_functions_0_ai1302_a110;
wire fp_functions_0_ai1302_a114_sumout;
wire fp_functions_0_ai1302_a115;
wire fp_functions_0_ai1302_a119_sumout;
wire fp_functions_0_ai1302_a120;
wire fp_functions_0_ai1302_a124_sumout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21_combout;
wire fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22_combout;
wire fp_functions_0_aMux_7_a2_combout;
wire fp_functions_0_aMux_6_a2_combout;
wire fp_functions_0_aMux_5_a2_combout;
wire fp_functions_0_aMux_4_a2_combout;
wire fp_functions_0_aMux_3_a2_combout;
wire fp_functions_0_aMux_2_a2_combout;
wire fp_functions_0_aMux_1_a2_combout;
wire fp_functions_0_aMux_0_a2_combout;
wire fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout;
wire fp_functions_0_ai1636_a0_combout;
wire fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0_combout;
wire fp_functions_0_ai1636_a1_combout;
wire fp_functions_0_ai1636_a2_combout;
wire fp_functions_0_ai1636_a3_combout;
wire fp_functions_0_ai1636_a4_combout;
wire fp_functions_0_ai1636_a5_combout;
wire fp_functions_0_ai1636_a6_combout;
wire fp_functions_0_ai1636_a7_combout;
wire fp_functions_0_ai1636_a8_combout;
wire fp_functions_0_ai1636_a9_combout;
wire fp_functions_0_ai1636_a10_combout;
wire fp_functions_0_ai1636_a11_combout;
wire fp_functions_0_ai1636_a12_combout;
wire fp_functions_0_ai1636_a13_combout;
wire fp_functions_0_ai1636_a14_combout;
wire fp_functions_0_ai1636_a15_combout;
wire fp_functions_0_ai1636_a16_combout;
wire fp_functions_0_ai1636_a17_combout;
wire fp_functions_0_ai1636_a18_combout;
wire fp_functions_0_ai1636_a19_combout;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq;
wire fp_functions_0_ai1636_a20_combout;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq;
wire fp_functions_0_ai1636_a21_combout;
wire fp_functions_0_ai1636_a22_combout;
wire fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0_combout;
wire fp_functions_0_aadd_2_a0_combout;
wire fp_functions_0_aadd_2_a1_combout;
wire fp_functions_0_aadd_2_a2_combout;
wire fp_functions_0_aadd_2_a3_combout;
wire fp_functions_0_aadd_2_a4_combout;
wire fp_functions_0_aadd_2_a5_combout;
wire fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4_combout;
wire fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5_combout;
wire fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6_combout;
wire fp_functions_0_ai1207_a0_combout;
wire fp_functions_0_areduce_nor_3_acombout;
wire fp_functions_0_areduce_nor_4_acombout;
wire fp_functions_0_ai1636_a23_combout;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq;
wire fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq;
wire fp_functions_0_areduce_or_0_a0_combout;
wire fp_functions_0_areduce_or_0_a1_combout;
wire fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7_combout;
wire fp_functions_0_ai1302_a0_combout;
wire fp_functions_0_ai1302_a1_combout;
wire fp_functions_0_ai1208_a0_combout;
wire fp_functions_0_ai1040_a1_combout;
wire fp_functions_0_ai1039_a1_combout;
wire fp_functions_0_ai1038_a1_combout;
wire fp_functions_0_ai1041_a1_combout;
wire fp_functions_0_ai1041_a2_combout;
wire fp_functions_0_ai1041_a3_combout;
wire fp_functions_0_ai1037_a1_combout;
wire fp_functions_0_ai1040_a2_combout;
wire fp_functions_0_ai1039_a2_combout;
wire fp_functions_0_ai1037_a2_combout;
wire fp_functions_0_ai1044_a1_combout;
wire fp_functions_0_ai1042_a1_combout;
wire fp_functions_0_ai1043_a1_combout;
wire fp_functions_0_areduce_nor_2_acombout;
wire fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout;
wire fp_functions_0_ai1132_a0_combout;
wire fp_functions_0_ai1302_a2_combout;
wire fp_functions_0_ai1302_a3_combout;
wire fp_functions_0_ai1302_a4_combout;
wire fp_functions_0_ai1302_a5_combout;
wire fp_functions_0_ai1302_a6_combout;
wire fp_functions_0_ai1302_a7_combout;
wire fp_functions_0_ai1132_a1_combout;
wire fp_functions_0_ai1132_a2_combout;
wire fp_functions_0_ai1132_a3_combout;
wire fp_functions_0_ai1132_a4_combout;
wire fp_functions_0_ai1132_a5_combout;
wire fp_functions_0_ai1132_a6_combout;
wire fp_functions_0_ai1132_a7_combout;
wire fp_functions_0_ai1132_a8_combout;
wire fp_functions_0_ai1132_a9_combout;
wire fp_functions_0_ai1132_a10_combout;
wire fp_functions_0_ai1132_a11_combout;
wire fp_functions_0_ai1132_a12_combout;
wire fp_functions_0_ai1132_a13_combout;
wire fp_functions_0_ai1132_a14_combout;
wire fp_functions_0_ai1132_a15_combout;
wire fp_functions_0_ai1044_a2_combout;
wire fp_functions_0_areduce_nor_0_a0_combout;
wire fp_functions_0_areduce_nor_0_a1_combout;
wire fp_functions_0_areduce_nor_0_a2_combout;
wire fp_functions_0_areduce_nor_0_a3_combout;
wire fp_functions_0_areduce_nor_0_a4_combout;
wire fp_functions_0_areduce_nor_0_a5_combout;
wire fp_functions_0_areduce_nor_0_acombout;
wire fp_functions_0_ai904_a1_combout;
wire fp_functions_0_ai904_a2_combout;
wire fp_functions_0_ai906_a1_combout;
wire fp_functions_0_ai901_a1_combout;
wire fp_functions_0_ai901_a2_combout;
wire fp_functions_0_ai904_a3_combout;
wire fp_functions_0_ai908_a1_combout;
wire fp_functions_0_ai908_a2_combout;
wire fp_functions_0_ai900_a1_combout;
wire fp_functions_0_ai903_a1_combout;
wire fp_functions_0_ai902_a1_combout;
wire fp_functions_0_ai899_a1_combout;
wire fp_functions_0_ai899_a2_combout;
wire fp_functions_0_ai904_a4_combout;
wire fp_functions_0_ai904_a5_combout;
wire fp_functions_0_ai906_a2_combout;
wire fp_functions_0_ai906_a3_combout;
wire fp_functions_0_ai905_a1_combout;
wire fp_functions_0_ai903_a2_combout;
wire fp_functions_0_ai911_a1_combout;
wire fp_functions_0_ai910_a1_combout;
wire fp_functions_0_ai910_a2_combout;
wire fp_functions_0_ai909_a1_combout;
wire fp_functions_0_ai907_a1_combout;
wire fp_functions_0_ai912_a1_combout;
wire fp_functions_0_ai912_a2_combout;
wire fp_functions_0_ai913_a1_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0_combout;
wire fp_functions_0_areduce_nor_1_acombout;
wire fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14_combout;
wire fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15_combout;
wire fp_functions_0_ai914_a1_combout;
wire fp_functions_0_aadd_2_a5_wirecell_combout;
wire fp_functions_0_areduce_nor_3_a_wirecell_combout;
wire fp_functions_0_areduce_nor_4_a_wirecell_combout;


fourteennm_ff fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ainIsZero_uid12_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_4_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_4_a1.extended_lut = "off";
defparam fp_functions_0_aadd_4_a1.lut_mask = 64'h0000000000000000;
defparam fp_functions_0_aadd_4_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_5_a1.extended_lut = "off";
defparam fp_functions_0_aadd_5_a1.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_5_a1.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a151_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ainIsZero_uid12_fxpToFPTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_ainIsZero_uid12_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_ainIsZero_uid12_fxpToFPTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_ainIsZero_uid12_fxpToFPTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_3_a1(
	.dataa(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a157_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a1_sumout),
	.cout(fp_functions_0_aadd_3_a2),
	.shareout());
defparam fp_functions_0_aadd_3_a1.extended_lut = "off";
defparam fp_functions_0_aadd_3_a1.lut_mask = 64'h0000000000005555;
defparam fp_functions_0_aadd_3_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a7.extended_lut = "off";
defparam fp_functions_0_aadd_4_a7.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_4_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a7.extended_lut = "off";
defparam fp_functions_0_aadd_5_a7.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_5_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a6_sumout),
	.cout(fp_functions_0_aadd_3_a7),
	.shareout());
defparam fp_functions_0_aadd_3_a6.extended_lut = "off";
defparam fp_functions_0_aadd_3_a6.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a11_sumout),
	.cout(fp_functions_0_aadd_3_a12),
	.shareout());
defparam fp_functions_0_aadd_3_a11.extended_lut = "off";
defparam fp_functions_0_aadd_3_a11.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a16_sumout),
	.cout(fp_functions_0_aadd_3_a17),
	.shareout());
defparam fp_functions_0_aadd_3_a16.extended_lut = "off";
defparam fp_functions_0_aadd_3_a16.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a21_sumout),
	.cout(fp_functions_0_aadd_3_a22),
	.shareout());
defparam fp_functions_0_aadd_3_a21.extended_lut = "off";
defparam fp_functions_0_aadd_3_a21.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a26_sumout),
	.cout(fp_functions_0_aadd_3_a27),
	.shareout());
defparam fp_functions_0_aadd_3_a26.extended_lut = "off";
defparam fp_functions_0_aadd_3_a26.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a31_sumout),
	.cout(fp_functions_0_aadd_3_a32),
	.shareout());
defparam fp_functions_0_aadd_3_a31.extended_lut = "off";
defparam fp_functions_0_aadd_3_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a36_sumout),
	.cout(fp_functions_0_aadd_3_a37),
	.shareout());
defparam fp_functions_0_aadd_3_a36.extended_lut = "off";
defparam fp_functions_0_aadd_3_a36.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a41_sumout),
	.cout(fp_functions_0_aadd_3_a42),
	.shareout());
defparam fp_functions_0_aadd_3_a41.extended_lut = "off";
defparam fp_functions_0_aadd_3_a41.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a46_sumout),
	.cout(fp_functions_0_aadd_3_a47),
	.shareout());
defparam fp_functions_0_aadd_3_a46.extended_lut = "off";
defparam fp_functions_0_aadd_3_a46.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a51_sumout),
	.cout(fp_functions_0_aadd_3_a52),
	.shareout());
defparam fp_functions_0_aadd_3_a51.extended_lut = "off";
defparam fp_functions_0_aadd_3_a51.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a56_sumout),
	.cout(fp_functions_0_aadd_3_a57),
	.shareout());
defparam fp_functions_0_aadd_3_a56.extended_lut = "off";
defparam fp_functions_0_aadd_3_a56.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a61_sumout),
	.cout(fp_functions_0_aadd_3_a62),
	.shareout());
defparam fp_functions_0_aadd_3_a61.extended_lut = "off";
defparam fp_functions_0_aadd_3_a61.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a66_sumout),
	.cout(fp_functions_0_aadd_3_a67),
	.shareout());
defparam fp_functions_0_aadd_3_a66.extended_lut = "off";
defparam fp_functions_0_aadd_3_a66.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a71_sumout),
	.cout(fp_functions_0_aadd_3_a72),
	.shareout());
defparam fp_functions_0_aadd_3_a71.extended_lut = "off";
defparam fp_functions_0_aadd_3_a71.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a76_sumout),
	.cout(fp_functions_0_aadd_3_a77),
	.shareout());
defparam fp_functions_0_aadd_3_a76.extended_lut = "off";
defparam fp_functions_0_aadd_3_a76.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a81_sumout),
	.cout(fp_functions_0_aadd_3_a82),
	.shareout());
defparam fp_functions_0_aadd_3_a81.extended_lut = "off";
defparam fp_functions_0_aadd_3_a81.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a86_sumout),
	.cout(fp_functions_0_aadd_3_a87),
	.shareout());
defparam fp_functions_0_aadd_3_a86.extended_lut = "off";
defparam fp_functions_0_aadd_3_a86.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a91_sumout),
	.cout(fp_functions_0_aadd_3_a92),
	.shareout());
defparam fp_functions_0_aadd_3_a91.extended_lut = "off";
defparam fp_functions_0_aadd_3_a91.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a96_sumout),
	.cout(fp_functions_0_aadd_3_a97),
	.shareout());
defparam fp_functions_0_aadd_3_a96.extended_lut = "off";
defparam fp_functions_0_aadd_3_a96.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a101_sumout),
	.cout(fp_functions_0_aadd_3_a102),
	.shareout());
defparam fp_functions_0_aadd_3_a101.extended_lut = "off";
defparam fp_functions_0_aadd_3_a101.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a106_sumout),
	.cout(fp_functions_0_aadd_3_a107),
	.shareout());
defparam fp_functions_0_aadd_3_a106.extended_lut = "off";
defparam fp_functions_0_aadd_3_a106.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a111_sumout),
	.cout(fp_functions_0_aadd_3_a112),
	.shareout());
defparam fp_functions_0_aadd_3_a111.extended_lut = "off";
defparam fp_functions_0_aadd_3_a111.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a116_sumout),
	.cout(fp_functions_0_aadd_3_a117),
	.shareout());
defparam fp_functions_0_aadd_3_a116.extended_lut = "off";
defparam fp_functions_0_aadd_3_a116.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a116.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a121_sumout),
	.cout(fp_functions_0_aadd_3_a122),
	.shareout());
defparam fp_functions_0_aadd_3_a121.extended_lut = "off";
defparam fp_functions_0_aadd_3_a121.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a121.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a126_sumout),
	.cout(fp_functions_0_aadd_3_a127),
	.shareout());
defparam fp_functions_0_aadd_3_a126.extended_lut = "off";
defparam fp_functions_0_aadd_3_a126.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a126.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a131_sumout),
	.cout(fp_functions_0_aadd_3_a132),
	.shareout());
defparam fp_functions_0_aadd_3_a131.extended_lut = "off";
defparam fp_functions_0_aadd_3_a131.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a131.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a136_sumout),
	.cout(fp_functions_0_aadd_3_a137),
	.shareout());
defparam fp_functions_0_aadd_3_a136.extended_lut = "off";
defparam fp_functions_0_aadd_3_a136.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a136.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a141_sumout),
	.cout(fp_functions_0_aadd_3_a142),
	.shareout());
defparam fp_functions_0_aadd_3_a141.extended_lut = "off";
defparam fp_functions_0_aadd_3_a141.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a141.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a146_sumout),
	.cout(fp_functions_0_aadd_3_a147),
	.shareout());
defparam fp_functions_0_aadd_3_a146.extended_lut = "off";
defparam fp_functions_0_aadd_3_a146.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a146.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a151_sumout),
	.cout(fp_functions_0_aadd_3_a152),
	.shareout());
defparam fp_functions_0_aadd_3_a151.extended_lut = "off";
defparam fp_functions_0_aadd_3_a151.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a151.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a1_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq));
defparam fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_3_a157(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a157_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a157.extended_lut = "off";
defparam fp_functions_0_aadd_3_a157.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_3_a157.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a12.extended_lut = "off";
defparam fp_functions_0_aadd_4_a12.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_4_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a12.extended_lut = "off";
defparam fp_functions_0_aadd_5_a12.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a12.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a17_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a18_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a19_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a20_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a21_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a22_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a23_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a0_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a1_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a2_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a3_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a4_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a5_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a5_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a5_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a6_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a7_a_aq));
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPreRnd_uid14_fxpToFPTest_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a2_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_1_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_1_a0_a_aq));
defparam fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_1_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a(
	.clk(clk),
	.d(fp_functions_0_ai1207_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a59_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a124_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1636_a23_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_asticky_uid20_fxpToFPTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_or_0_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_asticky_uid20_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_asticky_uid20_fxpToFPTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_asticky_uid20_fxpToFPTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_3_a161_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_4_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a17.extended_lut = "off";
defparam fp_functions_0_aadd_4_a17.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_4_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a17.extended_lut = "off";
defparam fp_functions_0_aadd_5_a17.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a17.shared_arith = "off";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a119_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a54_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a114_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a49_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a109_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a44_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a104_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a39_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a99_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a34_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a94_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a29_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a89_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a24_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a84_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a19_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a79_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a14_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a74_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a(
	.clk(clk),
	.d(fp_functions_0_ai1208_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_4_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_3_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a_aq));
defparam fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a3_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_0_a0_a_aq));
defparam fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a(
	.clk(clk),
	.d(fp_functions_0_ai1038_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a(
	.clk(clk),
	.d(fp_functions_0_ai1041_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a(
	.clk(clk),
	.d(fp_functions_0_ai1040_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a(
	.clk(clk),
	.d(fp_functions_0_ai1039_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a(
	.clk(clk),
	.d(fp_functions_0_ai1037_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_ai1042_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_ai1043_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a64_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_3_a161(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a161_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_3_a161.extended_lut = "off";
defparam fp_functions_0_aadd_3_a161.lut_mask = 64'h0000000000000000;
defparam fp_functions_0_aadd_3_a161.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a22.extended_lut = "off";
defparam fp_functions_0_aadd_4_a22.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_4_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a22.extended_lut = "off";
defparam fp_functions_0_aadd_5_a22.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a22.shared_arith = "off";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai1132_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_ai1044_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_2_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_aq));
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_1_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_1_a0_a_aq));
defparam fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_1_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a4_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_0_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a(
	.clk(clk),
	.d(fp_functions_0_ai901_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai908_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a(
	.clk(clk),
	.d(fp_functions_0_ai900_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a(
	.clk(clk),
	.d(fp_functions_0_ai902_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a(
	.clk(clk),
	.d(fp_functions_0_ai899_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_ai904_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_ai906_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_ai905_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a(
	.clk(clk),
	.d(fp_functions_0_ai903_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai911_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai910_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai909_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai907_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai912_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai913_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq));
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_4_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a27.extended_lut = "off";
defparam fp_functions_0_aadd_4_a27.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_4_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a27.extended_lut = "off";
defparam fp_functions_0_aadd_5_a27.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a27.shared_arith = "off";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai914_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq));
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_1_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_0_a0_a_aq));
defparam fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a5_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a151_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a(
	.clk(clk),
	.d(fp_functions_0_aadd_0_a156_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a_aq));
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a_aq));
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_4_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a32.extended_lut = "off";
defparam fp_functions_0_aadd_4_a32.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_4_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a32.extended_lut = "off";
defparam fp_functions_0_aadd_5_a32.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a32.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a6_a_a0_a_aq));
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_0_a1(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[13]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a1_sumout),
	.cout(fp_functions_0_aadd_0_a2),
	.shareout());
defparam fp_functions_0_aadd_0_a1.extended_lut = "off";
defparam fp_functions_0_aadd_0_a1.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a6(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[19]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a6_sumout),
	.cout(fp_functions_0_aadd_0_a7),
	.shareout());
defparam fp_functions_0_aadd_0_a6.extended_lut = "off";
defparam fp_functions_0_aadd_0_a6.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a11(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[21]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a11_sumout),
	.cout(fp_functions_0_aadd_0_a12),
	.shareout());
defparam fp_functions_0_aadd_0_a11.extended_lut = "off";
defparam fp_functions_0_aadd_0_a11.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a16(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a16_sumout),
	.cout(fp_functions_0_aadd_0_a17),
	.shareout());
defparam fp_functions_0_aadd_0_a16.extended_lut = "off";
defparam fp_functions_0_aadd_0_a16.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a21(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[24]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a21_sumout),
	.cout(fp_functions_0_aadd_0_a22),
	.shareout());
defparam fp_functions_0_aadd_0_a21.extended_lut = "off";
defparam fp_functions_0_aadd_0_a21.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a26(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[23]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a26_sumout),
	.cout(fp_functions_0_aadd_0_a27),
	.shareout());
defparam fp_functions_0_aadd_0_a26.extended_lut = "off";
defparam fp_functions_0_aadd_0_a26.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a31(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a31_sumout),
	.cout(fp_functions_0_aadd_0_a32),
	.shareout());
defparam fp_functions_0_aadd_0_a31.extended_lut = "off";
defparam fp_functions_0_aadd_0_a31.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a36(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[20]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a36_sumout),
	.cout(fp_functions_0_aadd_0_a37),
	.shareout());
defparam fp_functions_0_aadd_0_a36.extended_lut = "off";
defparam fp_functions_0_aadd_0_a36.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a41(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a41_sumout),
	.cout(fp_functions_0_aadd_0_a42),
	.shareout());
defparam fp_functions_0_aadd_0_a41.extended_lut = "off";
defparam fp_functions_0_aadd_0_a41.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a46(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[15]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a46_sumout),
	.cout(fp_functions_0_aadd_0_a47),
	.shareout());
defparam fp_functions_0_aadd_0_a46.extended_lut = "off";
defparam fp_functions_0_aadd_0_a46.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a51(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[16]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a51_sumout),
	.cout(fp_functions_0_aadd_0_a52),
	.shareout());
defparam fp_functions_0_aadd_0_a51.extended_lut = "off";
defparam fp_functions_0_aadd_0_a51.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a56(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[11]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a56_sumout),
	.cout(fp_functions_0_aadd_0_a57),
	.shareout());
defparam fp_functions_0_aadd_0_a56.extended_lut = "off";
defparam fp_functions_0_aadd_0_a56.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a61(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[17]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a61_sumout),
	.cout(fp_functions_0_aadd_0_a62),
	.shareout());
defparam fp_functions_0_aadd_0_a61.extended_lut = "off";
defparam fp_functions_0_aadd_0_a61.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a66(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a66_sumout),
	.cout(fp_functions_0_aadd_0_a67),
	.shareout());
defparam fp_functions_0_aadd_0_a66.extended_lut = "off";
defparam fp_functions_0_aadd_0_a66.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a71(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a71_sumout),
	.cout(fp_functions_0_aadd_0_a72),
	.shareout());
defparam fp_functions_0_aadd_0_a71.extended_lut = "off";
defparam fp_functions_0_aadd_0_a71.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a76(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[12]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a76_sumout),
	.cout(fp_functions_0_aadd_0_a77),
	.shareout());
defparam fp_functions_0_aadd_0_a76.extended_lut = "off";
defparam fp_functions_0_aadd_0_a76.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a81(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[26]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a81_sumout),
	.cout(fp_functions_0_aadd_0_a82),
	.shareout());
defparam fp_functions_0_aadd_0_a81.extended_lut = "off";
defparam fp_functions_0_aadd_0_a81.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a86(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a86_sumout),
	.cout(fp_functions_0_aadd_0_a87),
	.shareout());
defparam fp_functions_0_aadd_0_a86.extended_lut = "off";
defparam fp_functions_0_aadd_0_a86.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a91(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a91_sumout),
	.cout(fp_functions_0_aadd_0_a92),
	.shareout());
defparam fp_functions_0_aadd_0_a91.extended_lut = "off";
defparam fp_functions_0_aadd_0_a91.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a96(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[0]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a96_sumout),
	.cout(fp_functions_0_aadd_0_a97),
	.shareout());
defparam fp_functions_0_aadd_0_a96.extended_lut = "off";
defparam fp_functions_0_aadd_0_a96.lut_mask = 64'h0000000050500F0F;
defparam fp_functions_0_aadd_0_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a101(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[3]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a101_sumout),
	.cout(fp_functions_0_aadd_0_a102),
	.shareout());
defparam fp_functions_0_aadd_0_a101.extended_lut = "off";
defparam fp_functions_0_aadd_0_a101.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a106(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a106_sumout),
	.cout(fp_functions_0_aadd_0_a107),
	.shareout());
defparam fp_functions_0_aadd_0_a106.extended_lut = "off";
defparam fp_functions_0_aadd_0_a106.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a111(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[7]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a111_sumout),
	.cout(fp_functions_0_aadd_0_a112),
	.shareout());
defparam fp_functions_0_aadd_0_a111.extended_lut = "off";
defparam fp_functions_0_aadd_0_a111.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a116(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[8]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a116_sumout),
	.cout(fp_functions_0_aadd_0_a117),
	.shareout());
defparam fp_functions_0_aadd_0_a116.extended_lut = "off";
defparam fp_functions_0_aadd_0_a116.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a116.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a121(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[9]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a121_sumout),
	.cout(fp_functions_0_aadd_0_a122),
	.shareout());
defparam fp_functions_0_aadd_0_a121.extended_lut = "off";
defparam fp_functions_0_aadd_0_a121.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a121.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a126(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a126_sumout),
	.cout(fp_functions_0_aadd_0_a127),
	.shareout());
defparam fp_functions_0_aadd_0_a126.extended_lut = "off";
defparam fp_functions_0_aadd_0_a126.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a126.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a131(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[5]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a131_sumout),
	.cout(fp_functions_0_aadd_0_a132),
	.shareout());
defparam fp_functions_0_aadd_0_a131.extended_lut = "off";
defparam fp_functions_0_aadd_0_a131.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a131.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a136_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_0_a136.extended_lut = "off";
defparam fp_functions_0_aadd_0_a136.lut_mask = 64'h0000000000000000;
defparam fp_functions_0_aadd_0_a136.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a141(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a141_sumout),
	.cout(fp_functions_0_aadd_0_a142),
	.shareout());
defparam fp_functions_0_aadd_0_a141.extended_lut = "off";
defparam fp_functions_0_aadd_0_a141.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a141.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a146(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[29]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a146_sumout),
	.cout(fp_functions_0_aadd_0_a147),
	.shareout());
defparam fp_functions_0_aadd_0_a146.extended_lut = "off";
defparam fp_functions_0_aadd_0_a146.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a146.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a151(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[28]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a157),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a151_sumout),
	.cout(fp_functions_0_aadd_0_a152),
	.shareout());
defparam fp_functions_0_aadd_0_a151.extended_lut = "off";
defparam fp_functions_0_aadd_0_a151.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a151.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a156(
	.dataa(!a[31]),
	.datab(gnd),
	.datac(!a[27]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a156_sumout),
	.cout(fp_functions_0_aadd_0_a157),
	.shareout());
defparam fp_functions_0_aadd_0_a156.extended_lut = "off";
defparam fp_functions_0_aadd_0_a156.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_0_a156.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a37.extended_lut = "off";
defparam fp_functions_0_aadd_4_a37.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_4_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a37.extended_lut = "off";
defparam fp_functions_0_aadd_5_a37.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a42.extended_lut = "off";
defparam fp_functions_0_aadd_4_a42.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_4_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a42.extended_lut = "off";
defparam fp_functions_0_aadd_5_a42.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_5_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_4_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_4_a47.extended_lut = "off";
defparam fp_functions_0_aadd_4_a47.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_4_a47.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_5_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_5_a47.extended_lut = "off";
defparam fp_functions_0_aadd_5_a47.lut_mask = 64'h00000000F0000FF0;
defparam fp_functions_0_aadd_5_a47.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a10(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_ai1302_a10_cout),
	.shareout());
defparam fp_functions_0_ai1302_a10.extended_lut = "off";
defparam fp_functions_0_ai1302_a10.lut_mask = 64'h0000000004150000;
defparam fp_functions_0_ai1302_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a14(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a10_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a14_sumout),
	.cout(fp_functions_0_ai1302_a15),
	.shareout());
defparam fp_functions_0_ai1302_a14.extended_lut = "off";
defparam fp_functions_0_ai1302_a14.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a19(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a15),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a19_sumout),
	.cout(fp_functions_0_ai1302_a20),
	.shareout());
defparam fp_functions_0_ai1302_a19.extended_lut = "off";
defparam fp_functions_0_ai1302_a19.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a24(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a20),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a24_sumout),
	.cout(fp_functions_0_ai1302_a25),
	.shareout());
defparam fp_functions_0_ai1302_a24.extended_lut = "off";
defparam fp_functions_0_ai1302_a24.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a24.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a29(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a25),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a29_sumout),
	.cout(fp_functions_0_ai1302_a30),
	.shareout());
defparam fp_functions_0_ai1302_a29.extended_lut = "off";
defparam fp_functions_0_ai1302_a29.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a29.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a34(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a30),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a34_sumout),
	.cout(fp_functions_0_ai1302_a35),
	.shareout());
defparam fp_functions_0_ai1302_a34.extended_lut = "off";
defparam fp_functions_0_ai1302_a34.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a34.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a39(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a35),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a39_sumout),
	.cout(fp_functions_0_ai1302_a40),
	.shareout());
defparam fp_functions_0_ai1302_a39.extended_lut = "off";
defparam fp_functions_0_ai1302_a39.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a39.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a44(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a40),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a44_sumout),
	.cout(fp_functions_0_ai1302_a45),
	.shareout());
defparam fp_functions_0_ai1302_a44.extended_lut = "off";
defparam fp_functions_0_ai1302_a44.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a44.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a49(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a45),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a49_sumout),
	.cout(fp_functions_0_ai1302_a50),
	.shareout());
defparam fp_functions_0_ai1302_a49.extended_lut = "off";
defparam fp_functions_0_ai1302_a49.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a49.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a54(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a50),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a54_sumout),
	.cout(fp_functions_0_ai1302_a55),
	.shareout());
defparam fp_functions_0_ai1302_a54.extended_lut = "off";
defparam fp_functions_0_ai1302_a54.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a54.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a59(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a55),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a59_sumout),
	.cout(fp_functions_0_ai1302_a60),
	.shareout());
defparam fp_functions_0_ai1302_a59.extended_lut = "off";
defparam fp_functions_0_ai1302_a59.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a59.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a64(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a60),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a64_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a64.extended_lut = "off";
defparam fp_functions_0_ai1302_a64.lut_mask = 64'h000000000000082A;
defparam fp_functions_0_ai1302_a64.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a70(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_ai1302_a70_cout),
	.shareout());
defparam fp_functions_0_ai1302_a70.extended_lut = "off";
defparam fp_functions_0_ai1302_a70.lut_mask = 64'h0000000004150000;
defparam fp_functions_0_ai1302_a70.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a74(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a70_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a74_sumout),
	.cout(fp_functions_0_ai1302_a75),
	.shareout());
defparam fp_functions_0_ai1302_a74.extended_lut = "off";
defparam fp_functions_0_ai1302_a74.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a74.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a79(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a75),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a79_sumout),
	.cout(fp_functions_0_ai1302_a80),
	.shareout());
defparam fp_functions_0_ai1302_a79.extended_lut = "off";
defparam fp_functions_0_ai1302_a79.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a79.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a84(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a80),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a84_sumout),
	.cout(fp_functions_0_ai1302_a85),
	.shareout());
defparam fp_functions_0_ai1302_a84.extended_lut = "off";
defparam fp_functions_0_ai1302_a84.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a84.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a89(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a85),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a89_sumout),
	.cout(fp_functions_0_ai1302_a90),
	.shareout());
defparam fp_functions_0_ai1302_a89.extended_lut = "off";
defparam fp_functions_0_ai1302_a89.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a89.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a94(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a90),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a94_sumout),
	.cout(fp_functions_0_ai1302_a95),
	.shareout());
defparam fp_functions_0_ai1302_a94.extended_lut = "off";
defparam fp_functions_0_ai1302_a94.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a94.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a99(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a95),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a99_sumout),
	.cout(fp_functions_0_ai1302_a100),
	.shareout());
defparam fp_functions_0_ai1302_a99.extended_lut = "off";
defparam fp_functions_0_ai1302_a99.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a99.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a104(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a100),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a104_sumout),
	.cout(fp_functions_0_ai1302_a105),
	.shareout());
defparam fp_functions_0_ai1302_a104.extended_lut = "off";
defparam fp_functions_0_ai1302_a104.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a104.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a109(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a105),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a109_sumout),
	.cout(fp_functions_0_ai1302_a110),
	.shareout());
defparam fp_functions_0_ai1302_a109.extended_lut = "off";
defparam fp_functions_0_ai1302_a109.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a109.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a114(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a110),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a114_sumout),
	.cout(fp_functions_0_ai1302_a115),
	.shareout());
defparam fp_functions_0_ai1302_a114.extended_lut = "off";
defparam fp_functions_0_ai1302_a114.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a114.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a119(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a115),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a119_sumout),
	.cout(fp_functions_0_ai1302_a120),
	.shareout());
defparam fp_functions_0_ai1302_a119.extended_lut = "off";
defparam fp_functions_0_ai1302_a119.lut_mask = 64'h000000000415082A;
defparam fp_functions_0_ai1302_a119.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a124(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_ai1302_a120),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_ai1302_a124_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a124.extended_lut = "off";
defparam fp_functions_0_ai1302_a124.lut_mask = 64'h000000000000082A;
defparam fp_functions_0_ai1302_a124.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a2_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a3_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a5_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a6_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a7_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a8_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a9_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a10_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a11_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a12_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a13_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a14_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a15_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a16_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a17_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a18_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a19_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a20_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a21_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22(
	.dataa(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_fracR_uid25_fxpToFPTest_b_1_q_a22_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22.extended_lut = "off";
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22.lut_mask = 64'h0020002000200020;
defparam fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_7_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_7_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_7_a2.extended_lut = "off";
defparam fp_functions_0_aMux_7_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_7_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_6_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a1_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_6_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_6_a2.extended_lut = "off";
defparam fp_functions_0_aMux_6_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_6_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_5_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a2_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_5_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_5_a2.extended_lut = "off";
defparam fp_functions_0_aMux_5_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_5_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_4_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a3_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_4_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_4_a2.extended_lut = "off";
defparam fp_functions_0_aMux_4_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_4_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_3_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a4_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_3_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_3_a2.extended_lut = "off";
defparam fp_functions_0_aMux_3_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_3_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a5_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a2.extended_lut = "off";
defparam fp_functions_0_aMux_2_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_2_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_1_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a6_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_1_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_1_a2.extended_lut = "off";
defparam fp_functions_0_aMux_1_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_1_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_0_a2(
	.dataa(!fp_functions_0_aredist6_expR_uid26_fxpToFPTest_b_1_q_a7_a_aq),
	.datab(!fp_functions_0_aredist8_inIsZero_uid12_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_4_a1_sumout),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_0_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_0_a2.extended_lut = "off";
defparam fp_functions_0_aMux_0_a2.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fp_functions_0_aMux_0_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0(
	.dataa(!areset),
	.datab(!en[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a0(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a0.extended_lut = "off";
defparam fp_functions_0_ai1636_a0.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_ai1636_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0(
	.dataa(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a1_a_aq),
	.datab(!fp_functions_0_aredist0_fracRnd_uid15_fxpToFPTest_merged_bit_select_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_asticky_uid20_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0.lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam fp_functions_0_aexpFracR_uid24_fxpToFPTest_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a1(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a1.extended_lut = "off";
defparam fp_functions_0_ai1636_a1.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a2(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a2.extended_lut = "off";
defparam fp_functions_0_ai1636_a2.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a3(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a3.extended_lut = "off";
defparam fp_functions_0_ai1636_a3.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a4(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a4.extended_lut = "off";
defparam fp_functions_0_ai1636_a4.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a5(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a5.extended_lut = "off";
defparam fp_functions_0_ai1636_a5.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a6(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a6.extended_lut = "off";
defparam fp_functions_0_ai1636_a6.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a7(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a7.extended_lut = "off";
defparam fp_functions_0_ai1636_a7.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a8(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a8.extended_lut = "off";
defparam fp_functions_0_ai1636_a8.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a9(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a9.extended_lut = "off";
defparam fp_functions_0_ai1636_a9.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a10(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a10.extended_lut = "off";
defparam fp_functions_0_ai1636_a10.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a11(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a11.extended_lut = "off";
defparam fp_functions_0_ai1636_a11.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a12(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a12.extended_lut = "off";
defparam fp_functions_0_ai1636_a12.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a13(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a13.extended_lut = "off";
defparam fp_functions_0_ai1636_a13.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a14(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a14.extended_lut = "off";
defparam fp_functions_0_ai1636_a14.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a15(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a15.extended_lut = "off";
defparam fp_functions_0_ai1636_a15.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a16(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a16.extended_lut = "off";
defparam fp_functions_0_ai1636_a16.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a17(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a17.extended_lut = "off";
defparam fp_functions_0_ai1636_a17.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a18(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a18.extended_lut = "off";
defparam fp_functions_0_ai1636_a18.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a19(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a19.extended_lut = "off";
defparam fp_functions_0_ai1636_a19.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a19.shared_arith = "off";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1636_a20(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a20.extended_lut = "off";
defparam fp_functions_0_ai1636_a20.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a20.shared_arith = "off";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_ai1636_a21(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a21.extended_lut = "off";
defparam fp_functions_0_ai1636_a21.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a22(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a22.extended_lut = "off";
defparam fp_functions_0_ai1636_a22.lut_mask = 64'h2727272727272727;
defparam fp_functions_0_ai1636_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_avCountFinal_uid86_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a0(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(!fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a0.extended_lut = "off";
defparam fp_functions_0_aadd_2_a0.lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam fp_functions_0_aadd_2_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a1(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(!fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq),
	.datad(!fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a1.extended_lut = "off";
defparam fp_functions_0_aadd_2_a1.lut_mask = 64'hF75DF75DF75DF75D;
defparam fp_functions_0_aadd_2_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a2(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(!fp_functions_0_aredist1_vCount_uid70_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq),
	.datad(!fp_functions_0_aredist2_vCount_uid63_lzcShifterZ1_uid10_fxpToFPTest_q_1_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a2.extended_lut = "off";
defparam fp_functions_0_aadd_2_a2.lut_mask = 64'h0008000800080008;
defparam fp_functions_0_aadd_2_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a3(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aadd_2_a2_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a3.extended_lut = "off";
defparam fp_functions_0_aadd_2_a3.lut_mask = 64'hD2D2D2D2D2D2D2D2;
defparam fp_functions_0_aadd_2_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a4(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a_aq),
	.datad(!fp_functions_0_aadd_2_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a4.extended_lut = "off";
defparam fp_functions_0_aadd_2_a4.lut_mask = 64'hF5D7F5D7F5D7F5D7;
defparam fp_functions_0_aadd_2_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a5(
	.dataa(!fp_functions_0_aredist5_vCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_q_4_q_a0_a_aq),
	.datab(!fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aredist4_vCount_uid49_lzcShifterZ1_uid10_fxpToFPTest_q_3_q_a0_a_aq),
	.datad(!fp_functions_0_aadd_2_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a5.extended_lut = "off";
defparam fp_functions_0_aadd_2_a5.lut_mask = 64'hAAA8AAA8AAA8AAA8;
defparam fp_functions_0_aadd_2_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4(
	.dataa(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datae(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4.extended_lut = "off";
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4.lut_mask = 64'hDFFF0000DFFF0000;
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5(
	.dataa(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datae(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5.extended_lut = "off";
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5.lut_mask = 64'hAAAA2AAAAAAA2AAA;
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6(
	.dataa(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datae(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6.extended_lut = "off";
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6.lut_mask = 64'hF0F070F0F0F070F0;
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1207_a0(
	.dataa(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4_combout),
	.datab(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5_combout),
	.datac(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1207_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1207_a0.extended_lut = "off";
defparam fp_functions_0_ai1207_a0.lut_mask = 64'hBABABABABABABABA;
defparam fp_functions_0_ai1207_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_3(
	.dataa(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_3_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_3.lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam fp_functions_0_areduce_nor_3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4(
	.dataa(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datae(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.dataf(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4.lut_mask = 64'h7555FFFFF555FFFF;
defparam fp_functions_0_areduce_nor_4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1636_a23(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1636_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1636_a23.extended_lut = "off";
defparam fp_functions_0_ai1636_a23.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_ai1636_a23.shared_arith = "off";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai1302_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fp_functions_0_aredist3_vCount_uid56_lzcShifterZ1_uid10_fxpToFPTest_q_2_delay_0_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq));
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_areduce_or_0_a0(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq),
	.datad(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_or_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_or_0_a0.extended_lut = "off";
defparam fp_functions_0_areduce_or_0_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_or_0_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_or_0_a1(
	.dataa(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datab(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq),
	.datac(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq),
	.datad(!fp_functions_0_avStagei_uid74_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq),
	.datae(!fp_functions_0_areduce_or_0_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_or_0_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_or_0_a1.extended_lut = "off";
defparam fp_functions_0_areduce_or_0_a1.lut_mask = 64'hFFFF1FFFFFFF1FFF;
defparam fp_functions_0_areduce_or_0_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7(
	.dataa(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datae(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7.extended_lut = "off";
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7.lut_mask = 64'hCCCC4CCCCCCC4CCC;
defparam fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7_combout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a0.extended_lut = "off";
defparam fp_functions_0_ai1302_a0.lut_mask = 64'h0A220A22AAAA0000;
defparam fp_functions_0_ai1302_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a1(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_a6_combout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a1.extended_lut = "off";
defparam fp_functions_0_ai1302_a1.lut_mask = 64'h0A220A22AAAA0000;
defparam fp_functions_0_ai1302_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1208_a0(
	.dataa(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_a4_combout),
	.datab(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_a5_combout),
	.datac(!fp_functions_0_avStagei_uid67_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_a7_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1208_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1208_a0.extended_lut = "off";
defparam fp_functions_0_ai1208_a0.lut_mask = 64'hDCDCDCDCDCDCDCDC;
defparam fp_functions_0_ai1208_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1040_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datad(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1040_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1040_a1.extended_lut = "off";
defparam fp_functions_0_ai1040_a1.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_ai1040_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1039_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(!fp_functions_0_ai1040_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1039_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1039_a1.extended_lut = "off";
defparam fp_functions_0_ai1039_a1.lut_mask = 64'h0808080808080808;
defparam fp_functions_0_ai1039_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1038_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datad(!fp_functions_0_ai1039_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1038_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1038_a1.extended_lut = "off";
defparam fp_functions_0_ai1038_a1.lut_mask = 64'h0F2F0F2F0F2F0F2F;
defparam fp_functions_0_ai1038_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1041_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datad(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1041_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1041_a1.extended_lut = "off";
defparam fp_functions_0_ai1041_a1.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_ai1041_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1041_a2(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datac(!fp_functions_0_ai1041_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1041_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1041_a2.extended_lut = "off";
defparam fp_functions_0_ai1041_a2.lut_mask = 64'h0808080808080808;
defparam fp_functions_0_ai1041_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1041_a3(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq),
	.datad(!fp_functions_0_ai1041_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1041_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1041_a3.extended_lut = "off";
defparam fp_functions_0_ai1041_a3.lut_mask = 64'h333B333B333B333B;
defparam fp_functions_0_ai1041_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1037_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datac(!fp_functions_0_ai1040_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1037_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1037_a1.extended_lut = "off";
defparam fp_functions_0_ai1037_a1.lut_mask = 64'h0808080808080808;
defparam fp_functions_0_ai1037_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1040_a2(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq),
	.datad(!fp_functions_0_ai1037_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1040_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1040_a2.extended_lut = "off";
defparam fp_functions_0_ai1040_a2.lut_mask = 64'h555D555D555D555D;
defparam fp_functions_0_ai1040_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1039_a2(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a29_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq),
	.datad(!fp_functions_0_ai1039_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1039_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1039_a2.extended_lut = "off";
defparam fp_functions_0_ai1039_a2.lut_mask = 64'h555D555D555D555D;
defparam fp_functions_0_ai1039_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1037_a2(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a28_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datad(!fp_functions_0_ai1037_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1037_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1037_a2.extended_lut = "off";
defparam fp_functions_0_ai1037_a2.lut_mask = 64'h333B333B333B333B;
defparam fp_functions_0_ai1037_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1044_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_ai1041_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1044_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1044_a1.extended_lut = "off";
defparam fp_functions_0_ai1044_a1.lut_mask = 64'h0808080808080808;
defparam fp_functions_0_ai1044_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1042_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq),
	.datad(!fp_functions_0_ai1044_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1042_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1042_a1.extended_lut = "off";
defparam fp_functions_0_ai1042_a1.lut_mask = 64'h555D555D555D555D;
defparam fp_functions_0_ai1042_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1043_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a25_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a27_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq),
	.datad(!fp_functions_0_ai1041_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1043_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1043_a1.extended_lut = "off";
defparam fp_functions_0_ai1043_a1.lut_mask = 64'h555D555D555D555D;
defparam fp_functions_0_ai1043_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_2(
	.dataa(!fp_functions_0_ai1040_a1_combout),
	.datab(!fp_functions_0_ai1041_a1_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_2_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_2.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_areduce_nor_2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_areduce_nor_2_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0.extended_lut = "off";
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a0(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a0.extended_lut = "off";
defparam fp_functions_0_ai1132_a0.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a2(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a2.extended_lut = "off";
defparam fp_functions_0_ai1302_a2.lut_mask = 64'h0000222200AA0A0A;
defparam fp_functions_0_ai1302_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a3(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a3.extended_lut = "off";
defparam fp_functions_0_ai1302_a3.lut_mask = 64'h000000AA22220A0A;
defparam fp_functions_0_ai1302_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a4(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a4.extended_lut = "off";
defparam fp_functions_0_ai1302_a4.lut_mask = 64'h002A002A002A002A;
defparam fp_functions_0_ai1302_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a5(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a30_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a31_a_aq),
	.datad(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a5.extended_lut = "off";
defparam fp_functions_0_ai1302_a5.lut_mask = 64'h002A002A002A002A;
defparam fp_functions_0_ai1302_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a6(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a6.extended_lut = "off";
defparam fp_functions_0_ai1302_a6.lut_mask = 64'h000A0022000A0022;
defparam fp_functions_0_ai1302_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1302_a7(
	.dataa(!areset),
	.datab(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.datac(!fp_functions_0_avStagei_uid60_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1302_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1302_a7.extended_lut = "off";
defparam fp_functions_0_ai1302_a7.lut_mask = 64'h0022000A0022000A;
defparam fp_functions_0_ai1302_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a1(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a1_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a1.extended_lut = "off";
defparam fp_functions_0_ai1132_a1.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a2(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a2.extended_lut = "off";
defparam fp_functions_0_ai1132_a2.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a3(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a3_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a3.extended_lut = "off";
defparam fp_functions_0_ai1132_a3.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a4(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a4_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a4.extended_lut = "off";
defparam fp_functions_0_ai1132_a4.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a5(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a5_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a5.extended_lut = "off";
defparam fp_functions_0_ai1132_a5.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a6(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a6_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a6.extended_lut = "off";
defparam fp_functions_0_ai1132_a6.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a7(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a7_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a7.extended_lut = "off";
defparam fp_functions_0_ai1132_a7.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a8(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a8_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a8.extended_lut = "off";
defparam fp_functions_0_ai1132_a8.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai1132_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a9(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a17_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a9_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a9.extended_lut = "off";
defparam fp_functions_0_ai1132_a9.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a10(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a18_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a10_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a10.extended_lut = "off";
defparam fp_functions_0_ai1132_a10.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a11(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a19_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a11_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a11.extended_lut = "off";
defparam fp_functions_0_ai1132_a11.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a12(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a20_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a12_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a12.extended_lut = "off";
defparam fp_functions_0_ai1132_a12.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a13(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a21_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a13_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a13.extended_lut = "off";
defparam fp_functions_0_ai1132_a13.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a14(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a22_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a14_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a14.extended_lut = "off";
defparam fp_functions_0_ai1132_a14.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1132_a15(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a23_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a15_a_aq),
	.datac(!fp_functions_0_areduce_nor_2_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1132_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1132_a15.extended_lut = "off";
defparam fp_functions_0_ai1132_a15.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai1132_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1044_a2(
	.dataa(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a26_a_aq),
	.datab(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a24_a_aq),
	.datac(!fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a16_a_aq),
	.datad(!fp_functions_0_ai1044_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1044_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1044_a2.extended_lut = "off";
defparam fp_functions_0_ai1044_a2.lut_mask = 64'h333B333B333B333B;
defparam fp_functions_0_ai1044_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a0(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a25_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a24_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a23_a_aq),
	.datad(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a22_a_aq),
	.datae(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a20_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_0_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a1(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a14_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a15_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a16_a_aq),
	.datad(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a11_a_aq),
	.datae(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a17_a_aq),
	.dataf(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a18_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a1.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_areduce_nor_0_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a2(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a2_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a3_a_aq),
	.datae(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a2.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_0_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a3(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a7_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a8_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a9_a_aq),
	.datad(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a10_a_aq),
	.datae(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a5_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a3.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_0_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a4(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a31_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a30_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a29_a_aq),
	.datad(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a28_a_aq),
	.datae(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a27_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a4.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_0_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a5(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a6_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a12_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a26_a_aq),
	.datad(!fp_functions_0_areduce_nor_0_a2_combout),
	.datae(!fp_functions_0_areduce_nor_0_a3_combout),
	.dataf(!fp_functions_0_areduce_nor_0_a4_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a5.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a5.lut_mask = 64'h0000000000000080;
defparam fp_functions_0_areduce_nor_0_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0(
	.dataa(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a13_a_aq),
	.datab(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a19_a_aq),
	.datac(!fp_functions_0_aredist9_y_uid9_fxpToFPTest_b_1_q_a21_a_aq),
	.datad(!fp_functions_0_areduce_nor_0_a0_combout),
	.datae(!fp_functions_0_areduce_nor_0_a1_combout),
	.dataf(!fp_functions_0_areduce_nor_0_a5_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0.lut_mask = 64'h0000000000000080;
defparam fp_functions_0_areduce_nor_0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai904_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a_aq),
	.datae(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai904_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai904_a1.extended_lut = "off";
defparam fp_functions_0_ai904_a1.lut_mask = 64'h2AAAAAAA2AAAAAAA;
defparam fp_functions_0_ai904_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai904_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a_aq),
	.datae(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai904_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai904_a2.extended_lut = "off";
defparam fp_functions_0_ai904_a2.lut_mask = 64'h2AAAAAAA2AAAAAAA;
defparam fp_functions_0_ai904_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai906_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a_aq),
	.datae(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai906_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai906_a1.extended_lut = "off";
defparam fp_functions_0_ai906_a1.lut_mask = 64'h2AAAAAAA2AAAAAAA;
defparam fp_functions_0_ai906_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai901_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a_aq),
	.datad(!fp_functions_0_ai904_a1_combout),
	.datae(!fp_functions_0_ai904_a2_combout),
	.dataf(!fp_functions_0_ai906_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai901_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai901_a1.extended_lut = "off";
defparam fp_functions_0_ai901_a1.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai901_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai901_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a_aq),
	.datae(!fp_functions_0_ai901_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai901_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai901_a2.extended_lut = "off";
defparam fp_functions_0_ai901_a2.lut_mask = 64'h00AA08AA00AA08AA;
defparam fp_functions_0_ai901_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai904_a3(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a_aq),
	.datae(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai904_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai904_a3.extended_lut = "off";
defparam fp_functions_0_ai904_a3.lut_mask = 64'h2AAAAAAA2AAAAAAA;
defparam fp_functions_0_ai904_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai908_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a_aq),
	.datad(!fp_functions_0_ai904_a1_combout),
	.datae(!fp_functions_0_ai906_a1_combout),
	.dataf(!fp_functions_0_ai904_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai908_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai908_a1.extended_lut = "off";
defparam fp_functions_0_ai908_a1.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai908_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai908_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a_aq),
	.datae(!fp_functions_0_ai908_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai908_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai908_a2.extended_lut = "off";
defparam fp_functions_0_ai908_a2.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai908_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai900_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a_aq),
	.datae(!fp_functions_0_ai901_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai900_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai900_a1.extended_lut = "off";
defparam fp_functions_0_ai900_a1.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai900_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai903_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a_aq),
	.datad(!fp_functions_0_ai904_a2_combout),
	.datae(!fp_functions_0_ai906_a1_combout),
	.dataf(!fp_functions_0_ai904_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai903_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai903_a1.extended_lut = "off";
defparam fp_functions_0_ai903_a1.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai903_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai902_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a_aq),
	.datae(!fp_functions_0_ai903_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai902_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai902_a1.extended_lut = "off";
defparam fp_functions_0_ai902_a1.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai902_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai899_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a30_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a29_a_aq),
	.datad(!fp_functions_0_ai904_a1_combout),
	.datae(!fp_functions_0_ai904_a2_combout),
	.dataf(!fp_functions_0_ai906_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai899_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai899_a1.extended_lut = "off";
defparam fp_functions_0_ai899_a1.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai899_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai899_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a_aq),
	.datae(!fp_functions_0_ai899_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai899_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai899_a2.extended_lut = "off";
defparam fp_functions_0_ai899_a2.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai899_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai904_a4(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a_aq),
	.datad(!fp_functions_0_ai904_a1_combout),
	.datae(!fp_functions_0_ai904_a2_combout),
	.dataf(!fp_functions_0_ai904_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai904_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai904_a4.extended_lut = "off";
defparam fp_functions_0_ai904_a4.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai904_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai904_a5(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a_aq),
	.datae(!fp_functions_0_ai904_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai904_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai904_a5.extended_lut = "off";
defparam fp_functions_0_ai904_a5.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai904_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai906_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a_aq),
	.datad(!fp_functions_0_ai904_a2_combout),
	.datae(!fp_functions_0_ai906_a1_combout),
	.dataf(!fp_functions_0_ai904_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai906_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai906_a2.extended_lut = "off";
defparam fp_functions_0_ai906_a2.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai906_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai906_a3(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a_aq),
	.datae(!fp_functions_0_ai906_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai906_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai906_a3.extended_lut = "off";
defparam fp_functions_0_ai906_a3.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai906_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai905_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a25_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a24_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a_aq),
	.datae(!fp_functions_0_ai906_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai905_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai905_a1.extended_lut = "off";
defparam fp_functions_0_ai905_a1.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai905_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai903_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a28_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a27_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a_aq),
	.datae(!fp_functions_0_ai903_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai903_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai903_a2.extended_lut = "off";
defparam fp_functions_0_ai903_a2.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai903_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai911_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a31_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a19_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a_aq),
	.datae(!fp_functions_0_ai899_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai911_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai911_a1.extended_lut = "off";
defparam fp_functions_0_ai911_a1.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai911_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai910_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a_aq),
	.datad(!fp_functions_0_ai904_a1_combout),
	.datae(!fp_functions_0_ai906_a1_combout),
	.dataf(!fp_functions_0_ai904_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai910_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai910_a1.extended_lut = "off";
defparam fp_functions_0_ai910_a1.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai910_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai910_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a_aq),
	.datae(!fp_functions_0_ai910_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai910_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai910_a2.extended_lut = "off";
defparam fp_functions_0_ai910_a2.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai910_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai909_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a21_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a20_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a_aq),
	.datae(!fp_functions_0_ai910_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai909_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai909_a1.extended_lut = "off";
defparam fp_functions_0_ai909_a1.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai909_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai907_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a23_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a22_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a_aq),
	.datae(!fp_functions_0_ai908_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai907_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai907_a1.extended_lut = "off";
defparam fp_functions_0_ai907_a1.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai907_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai912_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a_aq),
	.datad(!fp_functions_0_ai904_a1_combout),
	.datae(!fp_functions_0_ai904_a2_combout),
	.dataf(!fp_functions_0_ai904_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai912_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai912_a1.extended_lut = "off";
defparam fp_functions_0_ai912_a1.lut_mask = 64'hD500000000000000;
defparam fp_functions_0_ai912_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai912_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a_aq),
	.datae(!fp_functions_0_ai912_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai912_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai912_a2.extended_lut = "off";
defparam fp_functions_0_ai912_a2.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai912_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai913_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a18_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a17_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a_aq),
	.datae(!fp_functions_0_ai912_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai913_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai913_a1.extended_lut = "off";
defparam fp_functions_0_ai913_a1.lut_mask = 64'h0A0A0A8A0A0A0A8A;
defparam fp_functions_0_ai913_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1(
	.dataa(!fp_functions_0_ai904_a1_combout),
	.datab(!fp_functions_0_ai904_a2_combout),
	.datac(!fp_functions_0_ai906_a1_combout),
	.datad(!fp_functions_0_ai904_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_areduce_nor_1_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0.extended_lut = "off";
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0.lut_mask = 64'h7777777777777777;
defparam fp_functions_0_avStagei_uid53_lzcShifterZ1_uid10_fxpToFPTest_q_a2_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a6_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a4_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a8_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a1_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a5_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a3_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a7_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a9_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a10_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a11_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a12_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a13_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a14_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a15_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15.extended_lut = "off";
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_avStagei_uid46_lzcShifterZ1_uid10_fxpToFPTest_q_a0_a_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai914_a1(
	.dataa(!fp_functions_0_avCount_uid44_lzcShifterZ1_uid10_fxpToFPTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a16_a_aq),
	.datac(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a26_a_aq),
	.datad(!fp_functions_0_aredist10_y_uid9_fxpToFPTest_b_2_q_a0_a_aq),
	.datae(!fp_functions_0_ai904_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai914_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai914_a1.extended_lut = "off";
defparam fp_functions_0_ai914_a1.lut_mask = 64'h222222A2222222A2;
defparam fp_functions_0_ai914_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a5_wirecell(
	.dataa(!fp_functions_0_aadd_2_a5_combout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aadd_2_a5_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a5_wirecell.extended_lut = "off";
defparam fp_functions_0_aadd_2_a5_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fp_functions_0_aadd_2_a5_wirecell.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_3_a_wirecell(
	.dataa(!fp_functions_0_areduce_nor_3_acombout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_3_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_3_a_wirecell.extended_lut = "off";
defparam fp_functions_0_areduce_nor_3_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fp_functions_0_areduce_nor_3_a_wirecell.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4_a_wirecell(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4_a_wirecell.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fp_functions_0_areduce_nor_4_a_wirecell.shared_arith = "off";

assign q[30] = fp_functions_0_aMux_0_a2_combout;

assign q[29] = fp_functions_0_aMux_1_a2_combout;

assign q[28] = fp_functions_0_aMux_2_a2_combout;

assign q[27] = fp_functions_0_aMux_3_a2_combout;

assign q[26] = fp_functions_0_aMux_4_a2_combout;

assign q[25] = fp_functions_0_aMux_5_a2_combout;

assign q[24] = fp_functions_0_aMux_6_a2_combout;

assign q[23] = fp_functions_0_aMux_7_a2_combout;

assign q[0] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a0_combout;

assign q[10] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a10_combout;

assign q[11] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a11_combout;

assign q[12] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a12_combout;

assign q[13] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a13_combout;

assign q[14] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a14_combout;

assign q[15] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a15_combout;

assign q[16] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a16_combout;

assign q[17] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a17_combout;

assign q[18] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a18_combout;

assign q[19] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a19_combout;

assign q[1] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a1_combout;

assign q[20] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a20_combout;

assign q[21] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a21_combout;

assign q[22] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a22_combout;

assign q[2] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a2_combout;

assign q[3] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a3_combout;

assign q[4] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a4_combout;

assign q[5] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a5_combout;

assign q[6] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a6_combout;

assign q[7] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a7_combout;

assign q[8] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a8_combout;

assign q[9] = fp_functions_0_aoutRes_uid40_fxpToFPTest_q_a0_a_a9_combout;

assign q[31] = fp_functions_0_aredist11_signX_uid6_fxpToFPTest_b_7_adelay_signals_a0_a_a0_a_aq;

endmodule
